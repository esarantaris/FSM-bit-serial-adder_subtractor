* SPICE3 file created from inverter.ext - technology: scmos

.include ../usc-spice

M1000 out in Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=26p ps=22u 
M1001 out in GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=19p ps=18u 
C0 in gnd! 4.8fF

Vgnd1 GND 0 DC 0V
Vgnd2 gnd! 0 DC 0V
VVdd Vdd 0 DC 2.8V
Vin in 0 pulse(0 2.8 0ns 0.1ns 0.1ns 10ns 20ns)
.tran 5ns 40ns
.probe
.end

