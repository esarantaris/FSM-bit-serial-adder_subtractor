* SPICE3 file created from fullsub_isolator.ext - technology: scmos

M1000 SubB_0/SR2B_2/dff3B_7/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=14040p ps=11880u 
M1001 SubB_0/SR2B_2/dff3B_7/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=9348p ps=8856u 
M1002 SubB_0/SR2B_2/dff3B_7/gate_0/S SubB_0/SR2B_2/dff3B_7/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1003 SubB_0/SR2B_2/dff3B_7/gate_0/S SubB_0/SR2B_2/dff3B_7/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1004 SubB_0/SR2B_2/dff3B_7/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1005 SubB_0/SR2B_2/dff3B_7/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1006 SubB_0/SR2B_2/dff3B_7/gate_3/Gout SUM0 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1007 SubB_0/SR2B_2/dff3B_7/gate_3/Gout SUM0 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1008 SubB_0/SR2B_2/dff3B_7/gate_3/Gout fsm_0/CLK SubB_0/SR2B_2/dff3B_7/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1009 SubB_0/SR2B_2/dff3B_7/gate_3/Gout SubB_0/SR2B_2/dff3B_7/gate_1/S SubB_0/SR2B_2/dff3B_7/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1010 SubB_0/SR2B_2/dff3B_7/gate_2/Gout SubB_0/SR2B_2/dff3B_7/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1011 SubB_0/SR2B_2/dff3B_7/gate_2/Gout SubB_0/SR2B_2/dff3B_7/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1012 SubB_0/SR2B_2/dff3B_7/gate_2/Gout SubB_0/SR2B_2/dff3B_7/gate_2/S SubB_0/SR2B_2/dff3B_7/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1013 SubB_0/SR2B_2/dff3B_7/gate_2/Gout SubB_0/SR2B_2/dff3B_7/gate_0/S SubB_0/SR2B_2/dff3B_7/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1014 SubB_0/SR2B_2/dff3B_7/Qb SUM0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1015 SubB_0/SR2B_2/dff3B_7/Qb SUM0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1016 SUM0 SubB_0/SR2B_2/dff3B_7/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=124p pd=82u as=0p ps=0u 
M1017 SUM0 SubB_0/SR2B_2/dff3B_7/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=75p pd=66u as=0p ps=0u 
M1018 SubB_0/SR2B_2/dff3B_7/gate_3/Gin SubB_0/SR2B_2/dff3B_7/gate_1/S SubB_0/SR2B_2/dff3B_7/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1019 SubB_0/SR2B_2/dff3B_7/gate_3/Gin fsm_0/CLK SubB_0/SR2B_2/dff3B_7/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1020 SubB_0/SR2B_2/dff3B_7/gate_1/Gin SubB_0/SR2B_2/dff3B_7/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1021 SubB_0/SR2B_2/dff3B_7/gate_1/Gin SubB_0/SR2B_2/dff3B_7/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1022 SubB_0/SR2B_2/dff3B_7/gate_2/Gin SubB_0/SR2B_2/dff3B_7/gate_0/S SubB_0/SR2B_2/dff3B_7/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1023 SubB_0/SR2B_2/dff3B_7/gate_2/Gin SubB_0/SR2B_2/dff3B_7/gate_2/S SubB_0/SR2B_2/dff3B_7/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1024 SubB_0/SR2B_2/dff3B_7/gate_0/Gin SubB_0/SR2B_2/dff3B_7/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1025 SubB_0/SR2B_2/dff3B_7/gate_0/Gin SubB_0/SR2B_2/dff3B_7/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1026 SubB_0/SR2B_2/dff3B_7/inverter_11/in SubB_0/SR2B_2/dff3B_7/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1027 Vdd SubB_0/SR2B_2/dff3B_7/D SubB_0/SR2B_2/dff3B_7/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1028 SubB_0/SR2B_2/dff3B_7/nand2_0/a_n37_n6# SubB_0/SR2B_2/dff3B_7/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1029 SubB_0/SR2B_2/dff3B_7/inverter_11/in SubB_0/SR2B_2/dff3B_7/D SubB_0/SR2B_2/dff3B_7/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1030 SubB_0/SR2B_2/dff3B_7/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1031 SubB_0/SR2B_2/dff3B_7/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1032 SubB_0/SR2B_2/dff3B_6/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1033 SubB_0/SR2B_2/dff3B_6/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1034 SubB_0/SR2B_2/dff3B_6/gate_0/S SubB_0/SR2B_2/dff3B_6/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1035 SubB_0/SR2B_2/dff3B_6/gate_0/S SubB_0/SR2B_2/dff3B_6/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1036 SubB_0/SR2B_2/dff3B_6/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1037 SubB_0/SR2B_2/dff3B_6/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1038 SubB_0/SR2B_2/dff3B_6/gate_3/Gout SUM1 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1039 SubB_0/SR2B_2/dff3B_6/gate_3/Gout SUM1 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1040 SubB_0/SR2B_2/dff3B_6/gate_3/Gout fsm_0/CLK SubB_0/SR2B_2/dff3B_6/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1041 SubB_0/SR2B_2/dff3B_6/gate_3/Gout SubB_0/SR2B_2/dff3B_6/gate_1/S SubB_0/SR2B_2/dff3B_6/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1042 SubB_0/SR2B_2/dff3B_6/gate_2/Gout SubB_0/SR2B_2/dff3B_6/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1043 SubB_0/SR2B_2/dff3B_6/gate_2/Gout SubB_0/SR2B_2/dff3B_6/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1044 SubB_0/SR2B_2/dff3B_6/gate_2/Gout SubB_0/SR2B_2/dff3B_6/gate_2/S SubB_0/SR2B_2/dff3B_6/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1045 SubB_0/SR2B_2/dff3B_6/gate_2/Gout SubB_0/SR2B_2/dff3B_6/gate_0/S SubB_0/SR2B_2/dff3B_6/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1046 SubB_0/SR2B_2/dff3B_6/Qb SUM1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1047 SubB_0/SR2B_2/dff3B_6/Qb SUM1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1048 SUM1 SubB_0/SR2B_2/dff3B_6/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M1049 SUM1 SubB_0/SR2B_2/dff3B_6/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M1050 SubB_0/SR2B_2/dff3B_6/gate_3/Gin SubB_0/SR2B_2/dff3B_6/gate_1/S SubB_0/SR2B_2/dff3B_6/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1051 SubB_0/SR2B_2/dff3B_6/gate_3/Gin fsm_0/CLK SubB_0/SR2B_2/dff3B_6/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1052 SubB_0/SR2B_2/dff3B_6/gate_1/Gin SubB_0/SR2B_2/dff3B_6/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1053 SubB_0/SR2B_2/dff3B_6/gate_1/Gin SubB_0/SR2B_2/dff3B_6/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1054 SubB_0/SR2B_2/dff3B_6/gate_2/Gin SubB_0/SR2B_2/dff3B_6/gate_0/S SubB_0/SR2B_2/dff3B_6/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1055 SubB_0/SR2B_2/dff3B_6/gate_2/Gin SubB_0/SR2B_2/dff3B_6/gate_2/S SubB_0/SR2B_2/dff3B_6/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1056 SubB_0/SR2B_2/dff3B_6/gate_0/Gin SubB_0/SR2B_2/dff3B_6/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1057 SubB_0/SR2B_2/dff3B_6/gate_0/Gin SubB_0/SR2B_2/dff3B_6/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1058 SubB_0/SR2B_2/dff3B_6/inverter_11/in SubB_0/SR2B_2/dff3B_6/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1059 Vdd SubB_0/SR2B_2/dff3B_6/D SubB_0/SR2B_2/dff3B_6/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1060 SubB_0/SR2B_2/dff3B_6/nand2_0/a_n37_n6# SubB_0/SR2B_2/dff3B_6/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1061 SubB_0/SR2B_2/dff3B_6/inverter_11/in SubB_0/SR2B_2/dff3B_6/D SubB_0/SR2B_2/dff3B_6/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1062 SubB_0/SR2B_2/dff3B_6/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1063 SubB_0/SR2B_2/dff3B_6/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1064 SubB_0/SR2B_2/dff3B_5/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1065 SubB_0/SR2B_2/dff3B_5/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1066 SubB_0/SR2B_2/dff3B_5/gate_0/S SubB_0/SR2B_2/dff3B_5/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1067 SubB_0/SR2B_2/dff3B_5/gate_0/S SubB_0/SR2B_2/dff3B_5/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1068 SubB_0/SR2B_2/dff3B_5/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1069 SubB_0/SR2B_2/dff3B_5/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1070 SubB_0/SR2B_2/dff3B_5/gate_3/Gout SUM2 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1071 SubB_0/SR2B_2/dff3B_5/gate_3/Gout SUM2 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1072 SubB_0/SR2B_2/dff3B_5/gate_3/Gout fsm_0/CLK SubB_0/SR2B_2/dff3B_5/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1073 SubB_0/SR2B_2/dff3B_5/gate_3/Gout SubB_0/SR2B_2/dff3B_5/gate_1/S SubB_0/SR2B_2/dff3B_5/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1074 SubB_0/SR2B_2/dff3B_5/gate_2/Gout SubB_0/SR2B_2/dff3B_5/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1075 SubB_0/SR2B_2/dff3B_5/gate_2/Gout SubB_0/SR2B_2/dff3B_5/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1076 SubB_0/SR2B_2/dff3B_5/gate_2/Gout SubB_0/SR2B_2/dff3B_5/gate_2/S SubB_0/SR2B_2/dff3B_5/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1077 SubB_0/SR2B_2/dff3B_5/gate_2/Gout SubB_0/SR2B_2/dff3B_5/gate_0/S SubB_0/SR2B_2/dff3B_5/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1078 SubB_0/SR2B_2/dff3B_5/Qb SUM2 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1079 SubB_0/SR2B_2/dff3B_5/Qb SUM2 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1080 SUM2 SubB_0/SR2B_2/dff3B_5/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M1081 SUM2 SubB_0/SR2B_2/dff3B_5/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M1082 SubB_0/SR2B_2/dff3B_5/gate_3/Gin SubB_0/SR2B_2/dff3B_5/gate_1/S SubB_0/SR2B_2/dff3B_5/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1083 SubB_0/SR2B_2/dff3B_5/gate_3/Gin fsm_0/CLK SubB_0/SR2B_2/dff3B_5/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1084 SubB_0/SR2B_2/dff3B_5/gate_1/Gin SubB_0/SR2B_2/dff3B_5/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1085 SubB_0/SR2B_2/dff3B_5/gate_1/Gin SubB_0/SR2B_2/dff3B_5/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1086 SubB_0/SR2B_2/dff3B_5/gate_2/Gin SubB_0/SR2B_2/dff3B_5/gate_0/S SubB_0/SR2B_2/dff3B_5/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1087 SubB_0/SR2B_2/dff3B_5/gate_2/Gin SubB_0/SR2B_2/dff3B_5/gate_2/S SubB_0/SR2B_2/dff3B_5/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1088 SubB_0/SR2B_2/dff3B_5/gate_0/Gin SubB_0/SR2B_2/dff3B_5/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1089 SubB_0/SR2B_2/dff3B_5/gate_0/Gin SubB_0/SR2B_2/dff3B_5/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1090 SubB_0/SR2B_2/dff3B_5/inverter_11/in SubB_0/SR2B_2/dff3B_5/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1091 Vdd SubB_0/SR2B_2/dff3B_5/D SubB_0/SR2B_2/dff3B_5/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1092 SubB_0/SR2B_2/dff3B_5/nand2_0/a_n37_n6# SubB_0/SR2B_2/dff3B_5/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1093 SubB_0/SR2B_2/dff3B_5/inverter_11/in SubB_0/SR2B_2/dff3B_5/D SubB_0/SR2B_2/dff3B_5/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1094 SubB_0/SR2B_2/dff3B_5/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1095 SubB_0/SR2B_2/dff3B_5/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1096 SubB_0/SR2B_2/dff3B_4/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1097 SubB_0/SR2B_2/dff3B_4/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1098 SubB_0/SR2B_2/dff3B_4/gate_0/S SubB_0/SR2B_2/dff3B_4/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1099 SubB_0/SR2B_2/dff3B_4/gate_0/S SubB_0/SR2B_2/dff3B_4/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1100 SubB_0/SR2B_2/dff3B_4/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1101 SubB_0/SR2B_2/dff3B_4/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1102 SubB_0/SR2B_2/dff3B_4/gate_3/Gout SUM3 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1103 SubB_0/SR2B_2/dff3B_4/gate_3/Gout SUM3 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1104 SubB_0/SR2B_2/dff3B_4/gate_3/Gout fsm_0/CLK SubB_0/SR2B_2/dff3B_4/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1105 SubB_0/SR2B_2/dff3B_4/gate_3/Gout SubB_0/SR2B_2/dff3B_4/gate_1/S SubB_0/SR2B_2/dff3B_4/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1106 SubB_0/SR2B_2/dff3B_4/gate_2/Gout SubB_0/SR2B_2/dff3B_4/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1107 SubB_0/SR2B_2/dff3B_4/gate_2/Gout SubB_0/SR2B_2/dff3B_4/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1108 SubB_0/SR2B_2/dff3B_4/gate_2/Gout SubB_0/SR2B_2/dff3B_4/gate_2/S SubB_0/SR2B_2/dff3B_4/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1109 SubB_0/SR2B_2/dff3B_4/gate_2/Gout SubB_0/SR2B_2/dff3B_4/gate_0/S SubB_0/SR2B_2/dff3B_4/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1110 SubB_0/SR2B_2/dff3B_4/Qb SUM3 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1111 SubB_0/SR2B_2/dff3B_4/Qb SUM3 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1112 SUM3 SubB_0/SR2B_2/dff3B_4/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M1113 SUM3 SubB_0/SR2B_2/dff3B_4/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M1114 SubB_0/SR2B_2/dff3B_4/gate_3/Gin SubB_0/SR2B_2/dff3B_4/gate_1/S SubB_0/SR2B_2/dff3B_4/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1115 SubB_0/SR2B_2/dff3B_4/gate_3/Gin fsm_0/CLK SubB_0/SR2B_2/dff3B_4/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1116 SubB_0/SR2B_2/dff3B_4/gate_1/Gin SubB_0/SR2B_2/dff3B_4/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1117 SubB_0/SR2B_2/dff3B_4/gate_1/Gin SubB_0/SR2B_2/dff3B_4/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1118 SubB_0/SR2B_2/dff3B_4/gate_2/Gin SubB_0/SR2B_2/dff3B_4/gate_0/S SubB_0/SR2B_2/dff3B_4/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1119 SubB_0/SR2B_2/dff3B_4/gate_2/Gin SubB_0/SR2B_2/dff3B_4/gate_2/S SubB_0/SR2B_2/dff3B_4/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1120 SubB_0/SR2B_2/dff3B_4/gate_0/Gin SubB_0/SR2B_2/dff3B_4/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1121 SubB_0/SR2B_2/dff3B_4/gate_0/Gin SubB_0/SR2B_2/dff3B_4/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1122 SubB_0/SR2B_2/dff3B_4/inverter_11/in SubB_0/SR2B_2/dff3B_4/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1123 Vdd SubB_0/SR2B_2/dff3B_4/D SubB_0/SR2B_2/dff3B_4/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1124 SubB_0/SR2B_2/dff3B_4/nand2_0/a_n37_n6# SubB_0/SR2B_2/dff3B_4/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1125 SubB_0/SR2B_2/dff3B_4/inverter_11/in SubB_0/SR2B_2/dff3B_4/D SubB_0/SR2B_2/dff3B_4/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1126 SubB_0/SR2B_2/dff3B_4/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1127 SubB_0/SR2B_2/dff3B_4/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1128 SubB_0/SR2B_2/dff3B_3/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1129 SubB_0/SR2B_2/dff3B_3/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1130 SubB_0/SR2B_2/dff3B_3/gate_0/S SubB_0/SR2B_2/dff3B_3/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1131 SubB_0/SR2B_2/dff3B_3/gate_0/S SubB_0/SR2B_2/dff3B_3/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1132 SubB_0/SR2B_2/dff3B_3/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1133 SubB_0/SR2B_2/dff3B_3/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1134 SubB_0/SR2B_2/dff3B_3/gate_3/Gout SUM4 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1135 SubB_0/SR2B_2/dff3B_3/gate_3/Gout SUM4 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1136 SubB_0/SR2B_2/dff3B_3/gate_3/Gout fsm_0/CLK SubB_0/SR2B_2/dff3B_3/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1137 SubB_0/SR2B_2/dff3B_3/gate_3/Gout SubB_0/SR2B_2/dff3B_3/gate_1/S SubB_0/SR2B_2/dff3B_3/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1138 SubB_0/SR2B_2/dff3B_3/gate_2/Gout SubB_0/SR2B_2/dff3B_3/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1139 SubB_0/SR2B_2/dff3B_3/gate_2/Gout SubB_0/SR2B_2/dff3B_3/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1140 SubB_0/SR2B_2/dff3B_3/gate_2/Gout SubB_0/SR2B_2/dff3B_3/gate_2/S SubB_0/SR2B_2/dff3B_3/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1141 SubB_0/SR2B_2/dff3B_3/gate_2/Gout SubB_0/SR2B_2/dff3B_3/gate_0/S SubB_0/SR2B_2/dff3B_3/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1142 SubB_0/SR2B_2/dff3B_3/Qb SUM4 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1143 SubB_0/SR2B_2/dff3B_3/Qb SUM4 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1144 SUM4 SubB_0/SR2B_2/dff3B_3/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M1145 SUM4 SubB_0/SR2B_2/dff3B_3/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M1146 SubB_0/SR2B_2/dff3B_3/gate_3/Gin SubB_0/SR2B_2/dff3B_3/gate_1/S SubB_0/SR2B_2/dff3B_3/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1147 SubB_0/SR2B_2/dff3B_3/gate_3/Gin fsm_0/CLK SubB_0/SR2B_2/dff3B_3/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1148 SubB_0/SR2B_2/dff3B_3/gate_1/Gin SubB_0/SR2B_2/dff3B_3/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1149 SubB_0/SR2B_2/dff3B_3/gate_1/Gin SubB_0/SR2B_2/dff3B_3/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1150 SubB_0/SR2B_2/dff3B_3/gate_2/Gin SubB_0/SR2B_2/dff3B_3/gate_0/S SubB_0/SR2B_2/dff3B_3/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1151 SubB_0/SR2B_2/dff3B_3/gate_2/Gin SubB_0/SR2B_2/dff3B_3/gate_2/S SubB_0/SR2B_2/dff3B_3/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1152 SubB_0/SR2B_2/dff3B_3/gate_0/Gin SubB_0/SR2B_2/dff3B_3/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1153 SubB_0/SR2B_2/dff3B_3/gate_0/Gin SubB_0/SR2B_2/dff3B_3/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1154 SubB_0/SR2B_2/dff3B_3/inverter_11/in SubB_0/SR2B_2/dff3B_3/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1155 Vdd SubB_0/SR2B_2/dff3B_3/D SubB_0/SR2B_2/dff3B_3/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1156 SubB_0/SR2B_2/dff3B_3/nand2_0/a_n37_n6# SubB_0/SR2B_2/dff3B_3/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1157 SubB_0/SR2B_2/dff3B_3/inverter_11/in SubB_0/SR2B_2/dff3B_3/D SubB_0/SR2B_2/dff3B_3/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1158 SubB_0/SR2B_2/dff3B_3/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1159 SubB_0/SR2B_2/dff3B_3/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1160 SubB_0/SR2B_2/dff3B_2/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1161 SubB_0/SR2B_2/dff3B_2/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1162 SubB_0/SR2B_2/dff3B_2/gate_0/S SubB_0/SR2B_2/dff3B_2/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1163 SubB_0/SR2B_2/dff3B_2/gate_0/S SubB_0/SR2B_2/dff3B_2/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1164 SubB_0/SR2B_2/dff3B_2/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1165 SubB_0/SR2B_2/dff3B_2/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1166 SubB_0/SR2B_2/dff3B_2/gate_3/Gout SUM5 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1167 SubB_0/SR2B_2/dff3B_2/gate_3/Gout SUM5 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1168 SubB_0/SR2B_2/dff3B_2/gate_3/Gout fsm_0/CLK SubB_0/SR2B_2/dff3B_2/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1169 SubB_0/SR2B_2/dff3B_2/gate_3/Gout SubB_0/SR2B_2/dff3B_2/gate_1/S SubB_0/SR2B_2/dff3B_2/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1170 SubB_0/SR2B_2/dff3B_2/gate_2/Gout SubB_0/SR2B_2/dff3B_2/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1171 SubB_0/SR2B_2/dff3B_2/gate_2/Gout SubB_0/SR2B_2/dff3B_2/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1172 SubB_0/SR2B_2/dff3B_2/gate_2/Gout SubB_0/SR2B_2/dff3B_2/gate_2/S SubB_0/SR2B_2/dff3B_2/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1173 SubB_0/SR2B_2/dff3B_2/gate_2/Gout SubB_0/SR2B_2/dff3B_2/gate_0/S SubB_0/SR2B_2/dff3B_2/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1174 SubB_0/SR2B_2/dff3B_2/Qb SUM5 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1175 SubB_0/SR2B_2/dff3B_2/Qb SUM5 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1176 SUM5 SubB_0/SR2B_2/dff3B_2/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M1177 SUM5 SubB_0/SR2B_2/dff3B_2/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M1178 SubB_0/SR2B_2/dff3B_2/gate_3/Gin SubB_0/SR2B_2/dff3B_2/gate_1/S SubB_0/SR2B_2/dff3B_2/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1179 SubB_0/SR2B_2/dff3B_2/gate_3/Gin fsm_0/CLK SubB_0/SR2B_2/dff3B_2/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1180 SubB_0/SR2B_2/dff3B_2/gate_1/Gin SubB_0/SR2B_2/dff3B_2/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1181 SubB_0/SR2B_2/dff3B_2/gate_1/Gin SubB_0/SR2B_2/dff3B_2/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1182 SubB_0/SR2B_2/dff3B_2/gate_2/Gin SubB_0/SR2B_2/dff3B_2/gate_0/S SubB_0/SR2B_2/dff3B_2/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1183 SubB_0/SR2B_2/dff3B_2/gate_2/Gin SubB_0/SR2B_2/dff3B_2/gate_2/S SubB_0/SR2B_2/dff3B_2/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1184 SubB_0/SR2B_2/dff3B_2/gate_0/Gin SubB_0/SR2B_2/dff3B_2/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1185 SubB_0/SR2B_2/dff3B_2/gate_0/Gin SubB_0/SR2B_2/dff3B_2/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1186 SubB_0/SR2B_2/dff3B_2/inverter_11/in SubB_0/SR2B_2/dff3B_2/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1187 Vdd SubB_0/SR2B_2/dff3B_2/D SubB_0/SR2B_2/dff3B_2/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1188 SubB_0/SR2B_2/dff3B_2/nand2_0/a_n37_n6# SubB_0/SR2B_2/dff3B_2/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1189 SubB_0/SR2B_2/dff3B_2/inverter_11/in SubB_0/SR2B_2/dff3B_2/D SubB_0/SR2B_2/dff3B_2/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1190 SubB_0/SR2B_2/dff3B_2/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1191 SubB_0/SR2B_2/dff3B_2/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1192 SubB_0/SR2B_2/dff3B_1/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1193 SubB_0/SR2B_2/dff3B_1/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1194 SubB_0/SR2B_2/dff3B_1/gate_0/S SubB_0/SR2B_2/dff3B_1/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1195 SubB_0/SR2B_2/dff3B_1/gate_0/S SubB_0/SR2B_2/dff3B_1/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1196 SubB_0/SR2B_2/dff3B_1/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1197 SubB_0/SR2B_2/dff3B_1/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1198 SubB_0/SR2B_2/dff3B_1/gate_3/Gout SUM6 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1199 SubB_0/SR2B_2/dff3B_1/gate_3/Gout SUM6 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1200 SubB_0/SR2B_2/dff3B_1/gate_3/Gout fsm_0/CLK SubB_0/SR2B_2/dff3B_1/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1201 SubB_0/SR2B_2/dff3B_1/gate_3/Gout SubB_0/SR2B_2/dff3B_1/gate_1/S SubB_0/SR2B_2/dff3B_1/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1202 SubB_0/SR2B_2/dff3B_1/gate_2/Gout SubB_0/SR2B_2/dff3B_1/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1203 SubB_0/SR2B_2/dff3B_1/gate_2/Gout SubB_0/SR2B_2/dff3B_1/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1204 SubB_0/SR2B_2/dff3B_1/gate_2/Gout SubB_0/SR2B_2/dff3B_1/gate_2/S SubB_0/SR2B_2/dff3B_1/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1205 SubB_0/SR2B_2/dff3B_1/gate_2/Gout SubB_0/SR2B_2/dff3B_1/gate_0/S SubB_0/SR2B_2/dff3B_1/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1206 SubB_0/SR2B_2/dff3B_1/Qb SUM6 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1207 SubB_0/SR2B_2/dff3B_1/Qb SUM6 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1208 SUM6 SubB_0/SR2B_2/dff3B_1/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M1209 SUM6 SubB_0/SR2B_2/dff3B_1/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M1210 SubB_0/SR2B_2/dff3B_1/gate_3/Gin SubB_0/SR2B_2/dff3B_1/gate_1/S SubB_0/SR2B_2/dff3B_1/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1211 SubB_0/SR2B_2/dff3B_1/gate_3/Gin fsm_0/CLK SubB_0/SR2B_2/dff3B_1/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1212 SubB_0/SR2B_2/dff3B_1/gate_1/Gin SubB_0/SR2B_2/dff3B_1/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1213 SubB_0/SR2B_2/dff3B_1/gate_1/Gin SubB_0/SR2B_2/dff3B_1/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1214 SubB_0/SR2B_2/dff3B_1/gate_2/Gin SubB_0/SR2B_2/dff3B_1/gate_0/S SubB_0/SR2B_2/dff3B_1/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1215 SubB_0/SR2B_2/dff3B_1/gate_2/Gin SubB_0/SR2B_2/dff3B_1/gate_2/S SubB_0/SR2B_2/dff3B_1/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1216 SubB_0/SR2B_2/dff3B_1/gate_0/Gin SubB_0/SR2B_2/dff3B_1/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1217 SubB_0/SR2B_2/dff3B_1/gate_0/Gin SubB_0/SR2B_2/dff3B_1/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1218 SubB_0/SR2B_2/dff3B_1/inverter_11/in SubB_0/SR2B_2/dff3B_1/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1219 Vdd SubB_0/SR2B_2/dff3B_1/D SubB_0/SR2B_2/dff3B_1/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1220 SubB_0/SR2B_2/dff3B_1/nand2_0/a_n37_n6# SubB_0/SR2B_2/dff3B_1/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1221 SubB_0/SR2B_2/dff3B_1/inverter_11/in SubB_0/SR2B_2/dff3B_1/D SubB_0/SR2B_2/dff3B_1/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1222 SubB_0/SR2B_2/dff3B_1/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1223 SubB_0/SR2B_2/dff3B_1/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1224 SubB_0/SR2B_2/dff3B_0/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1225 SubB_0/SR2B_2/dff3B_0/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1226 SubB_0/SR2B_2/dff3B_0/gate_0/S SubB_0/SR2B_2/dff3B_0/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1227 SubB_0/SR2B_2/dff3B_0/gate_0/S SubB_0/SR2B_2/dff3B_0/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1228 SubB_0/SR2B_2/dff3B_0/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1229 SubB_0/SR2B_2/dff3B_0/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1230 SubB_0/SR2B_2/dff3B_0/gate_3/Gout SUM7 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1231 SubB_0/SR2B_2/dff3B_0/gate_3/Gout SUM7 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1232 SubB_0/SR2B_2/dff3B_0/gate_3/Gout fsm_0/CLK SubB_0/SR2B_2/dff3B_0/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1233 SubB_0/SR2B_2/dff3B_0/gate_3/Gout SubB_0/SR2B_2/dff3B_0/gate_1/S SubB_0/SR2B_2/dff3B_0/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1234 SubB_0/SR2B_2/dff3B_0/gate_2/Gout SubB_0/SR2B_2/dff3B_0/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1235 SubB_0/SR2B_2/dff3B_0/gate_2/Gout SubB_0/SR2B_2/dff3B_0/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1236 SubB_0/SR2B_2/dff3B_0/gate_2/Gout SubB_0/SR2B_2/dff3B_0/gate_2/S SubB_0/SR2B_2/dff3B_0/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1237 SubB_0/SR2B_2/dff3B_0/gate_2/Gout SubB_0/SR2B_2/dff3B_0/gate_0/S SubB_0/SR2B_2/dff3B_0/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1238 SubB_0/SR2B_2/dff3B_0/Qb SUM7 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1239 SubB_0/SR2B_2/dff3B_0/Qb SUM7 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1240 SUM7 SubB_0/SR2B_2/dff3B_0/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=124p pd=82u as=0p ps=0u 
M1241 SUM7 SubB_0/SR2B_2/dff3B_0/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=75p pd=66u as=0p ps=0u 
M1242 SubB_0/SR2B_2/dff3B_0/gate_3/Gin SubB_0/SR2B_2/dff3B_0/gate_1/S SubB_0/SR2B_2/dff3B_0/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1243 SubB_0/SR2B_2/dff3B_0/gate_3/Gin fsm_0/CLK SubB_0/SR2B_2/dff3B_0/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1244 SubB_0/SR2B_2/dff3B_0/gate_1/Gin SubB_0/SR2B_2/dff3B_0/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1245 SubB_0/SR2B_2/dff3B_0/gate_1/Gin SubB_0/SR2B_2/dff3B_0/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1246 SubB_0/SR2B_2/dff3B_0/gate_2/Gin SubB_0/SR2B_2/dff3B_0/gate_0/S SubB_0/SR2B_2/dff3B_0/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1247 SubB_0/SR2B_2/dff3B_0/gate_2/Gin SubB_0/SR2B_2/dff3B_0/gate_2/S SubB_0/SR2B_2/dff3B_0/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1248 SubB_0/SR2B_2/dff3B_0/gate_0/Gin SubB_0/SR2B_2/dff3B_0/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1249 SubB_0/SR2B_2/dff3B_0/gate_0/Gin SubB_0/SR2B_2/dff3B_0/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1250 SubB_0/SR2B_2/dff3B_0/inverter_11/in SubB_0/SR2B_2/dff3B_0/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1251 Vdd SubB_0/SR2B_2/dff3B_0/D SubB_0/SR2B_2/dff3B_0/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1252 SubB_0/SR2B_2/dff3B_0/nand2_0/a_n37_n6# SubB_0/SR2B_2/dff3B_0/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1253 SubB_0/SR2B_2/dff3B_0/inverter_11/in SubB_0/SR2B_2/dff3B_0/D SubB_0/SR2B_2/dff3B_0/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1254 SubB_0/SR2B_2/dff3B_0/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1255 SubB_0/SR2B_2/dff3B_0/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1256 SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Min2 nor2_0/out SUM0 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M1257 SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Min2 SubB_0/SR2B_2/mux4x1_7/mux2x1_1/Smb SUM0 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M1258 SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Min2 SubB_0/SR2B_2/mux4x1_7/mux2x1_1/Smb SL Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M1259 SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Min2 nor2_0/out SL Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M1260 SubB_0/SR2B_2/dff3B_7/D SS0 SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M1261 SubB_0/SR2B_2/dff3B_7/D SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Smb SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M1262 SubB_0/SR2B_2/dff3B_7/D SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Smb SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M1263 SubB_0/SR2B_2/dff3B_7/D SS0 SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M1264 SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Min1 nor2_0/out SUM1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1265 SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Min1 SubB_0/SR2B_2/mux4x1_7/mux2x1_1/Smb SUM1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1266 SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Min1 SubB_0/SR2B_2/mux4x1_7/mux2x1_1/Smb D7 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M1267 SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Min1 nor2_0/out D7 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M1268 SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Smb SS0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1269 SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Smb SS0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1270 SubB_0/SR2B_2/mux4x1_7/mux2x1_1/Smb nor2_0/out Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1271 SubB_0/SR2B_2/mux4x1_7/mux2x1_1/Smb nor2_0/out GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1272 SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Min2 nor2_0/out SUM1 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M1273 SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Min2 SubB_0/SR2B_2/mux4x1_6/mux2x1_1/Smb SUM1 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M1274 SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Min2 SubB_0/SR2B_2/mux4x1_6/mux2x1_1/Smb SUM0 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1275 SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Min2 nor2_0/out SUM0 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1276 SubB_0/SR2B_2/dff3B_6/D SS0 SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M1277 SubB_0/SR2B_2/dff3B_6/D SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Smb SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M1278 SubB_0/SR2B_2/dff3B_6/D SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Smb SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M1279 SubB_0/SR2B_2/dff3B_6/D SS0 SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M1280 SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Min1 nor2_0/out SUM2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1281 SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Min1 SubB_0/SR2B_2/mux4x1_6/mux2x1_1/Smb SUM2 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1282 SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Min1 SubB_0/SR2B_2/mux4x1_6/mux2x1_1/Smb D6 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M1283 SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Min1 nor2_0/out D6 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M1284 SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Smb SS0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1285 SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Smb SS0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1286 SubB_0/SR2B_2/mux4x1_6/mux2x1_1/Smb nor2_0/out Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1287 SubB_0/SR2B_2/mux4x1_6/mux2x1_1/Smb nor2_0/out GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1288 SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Min2 nor2_0/out SUM2 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M1289 SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Min2 SubB_0/SR2B_2/mux4x1_5/mux2x1_1/Smb SUM2 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M1290 SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Min2 SubB_0/SR2B_2/mux4x1_5/mux2x1_1/Smb SUM1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1291 SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Min2 nor2_0/out SUM1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1292 SubB_0/SR2B_2/dff3B_5/D SS0 SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M1293 SubB_0/SR2B_2/dff3B_5/D SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Smb SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M1294 SubB_0/SR2B_2/dff3B_5/D SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Smb SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M1295 SubB_0/SR2B_2/dff3B_5/D SS0 SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M1296 SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Min1 nor2_0/out SUM3 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1297 SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Min1 SubB_0/SR2B_2/mux4x1_5/mux2x1_1/Smb SUM3 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1298 SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Min1 SubB_0/SR2B_2/mux4x1_5/mux2x1_1/Smb D5 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M1299 SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Min1 nor2_0/out D5 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M1300 SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Smb SS0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1301 SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Smb SS0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1302 SubB_0/SR2B_2/mux4x1_5/mux2x1_1/Smb nor2_0/out Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1303 SubB_0/SR2B_2/mux4x1_5/mux2x1_1/Smb nor2_0/out GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1304 SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Min2 nor2_0/out SUM3 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M1305 SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Min2 SubB_0/SR2B_2/mux4x1_4/mux2x1_1/Smb SUM3 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M1306 SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Min2 SubB_0/SR2B_2/mux4x1_4/mux2x1_1/Smb SUM2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1307 SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Min2 nor2_0/out SUM2 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1308 SubB_0/SR2B_2/dff3B_4/D SS0 SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M1309 SubB_0/SR2B_2/dff3B_4/D SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Smb SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M1310 SubB_0/SR2B_2/dff3B_4/D SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Smb SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M1311 SubB_0/SR2B_2/dff3B_4/D SS0 SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M1312 SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Min1 nor2_0/out SUM4 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1313 SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Min1 SubB_0/SR2B_2/mux4x1_4/mux2x1_1/Smb SUM4 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1314 SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Min1 SubB_0/SR2B_2/mux4x1_4/mux2x1_1/Smb D4 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M1315 SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Min1 nor2_0/out D4 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M1316 SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Smb SS0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1317 SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Smb SS0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1318 SubB_0/SR2B_2/mux4x1_4/mux2x1_1/Smb nor2_0/out Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1319 SubB_0/SR2B_2/mux4x1_4/mux2x1_1/Smb nor2_0/out GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1320 SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Min2 nor2_0/out SUM4 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M1321 SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Min2 SubB_0/SR2B_2/mux4x1_3/mux2x1_1/Smb SUM4 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M1322 SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Min2 SubB_0/SR2B_2/mux4x1_3/mux2x1_1/Smb SUM3 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1323 SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Min2 nor2_0/out SUM3 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1324 SubB_0/SR2B_2/dff3B_3/D SS0 SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M1325 SubB_0/SR2B_2/dff3B_3/D SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Smb SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M1326 SubB_0/SR2B_2/dff3B_3/D SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Smb SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M1327 SubB_0/SR2B_2/dff3B_3/D SS0 SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M1328 SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Min1 nor2_0/out SUM5 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1329 SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Min1 SubB_0/SR2B_2/mux4x1_3/mux2x1_1/Smb SUM5 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1330 SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Min1 SubB_0/SR2B_2/mux4x1_3/mux2x1_1/Smb D3 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M1331 SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Min1 nor2_0/out D3 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M1332 SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Smb SS0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1333 SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Smb SS0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1334 SubB_0/SR2B_2/mux4x1_3/mux2x1_1/Smb nor2_0/out Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1335 SubB_0/SR2B_2/mux4x1_3/mux2x1_1/Smb nor2_0/out GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1336 SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Min2 nor2_0/out SUM5 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M1337 SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Min2 SubB_0/SR2B_2/mux4x1_2/mux2x1_1/Smb SUM5 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M1338 SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Min2 SubB_0/SR2B_2/mux4x1_2/mux2x1_1/Smb SUM4 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1339 SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Min2 nor2_0/out SUM4 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1340 SubB_0/SR2B_2/dff3B_2/D SS0 SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M1341 SubB_0/SR2B_2/dff3B_2/D SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Smb SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M1342 SubB_0/SR2B_2/dff3B_2/D SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Smb SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M1343 SubB_0/SR2B_2/dff3B_2/D SS0 SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M1344 SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Min1 nor2_0/out SUM6 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1345 SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Min1 SubB_0/SR2B_2/mux4x1_2/mux2x1_1/Smb SUM6 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1346 SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Min1 SubB_0/SR2B_2/mux4x1_2/mux2x1_1/Smb D2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M1347 SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Min1 nor2_0/out D2 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M1348 SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Smb SS0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1349 SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Smb SS0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1350 SubB_0/SR2B_2/mux4x1_2/mux2x1_1/Smb nor2_0/out Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1351 SubB_0/SR2B_2/mux4x1_2/mux2x1_1/Smb nor2_0/out GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1352 SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Min2 nor2_0/out SUM6 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M1353 SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Min2 SubB_0/SR2B_2/mux4x1_1/mux2x1_1/Smb SUM6 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M1354 SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Min2 SubB_0/SR2B_2/mux4x1_1/mux2x1_1/Smb SUM5 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1355 SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Min2 nor2_0/out SUM5 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1356 SubB_0/SR2B_2/dff3B_1/D SS0 SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M1357 SubB_0/SR2B_2/dff3B_1/D SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Smb SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M1358 SubB_0/SR2B_2/dff3B_1/D SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Smb SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M1359 SubB_0/SR2B_2/dff3B_1/D SS0 SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M1360 SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Min1 nor2_0/out SUM7 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1361 SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Min1 SubB_0/SR2B_2/mux4x1_1/mux2x1_1/Smb SUM7 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1362 SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Min1 SubB_0/SR2B_2/mux4x1_1/mux2x1_1/Smb D1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M1363 SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Min1 nor2_0/out D1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M1364 SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Smb SS0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1365 SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Smb SS0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1366 SubB_0/SR2B_2/mux4x1_1/mux2x1_1/Smb nor2_0/out Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1367 SubB_0/SR2B_2/mux4x1_1/mux2x1_1/Smb nor2_0/out GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1368 SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Min2 nor2_0/out SUM7 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M1369 SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Min2 SubB_0/SR2B_2/mux4x1_0/mux2x1_1/Smb SUM7 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M1370 SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Min2 SubB_0/SR2B_2/mux4x1_0/mux2x1_1/Smb SUM6 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1371 SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Min2 nor2_0/out SUM6 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1372 SubB_0/SR2B_2/dff3B_0/D SS0 SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M1373 SubB_0/SR2B_2/dff3B_0/D SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Smb SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M1374 SubB_0/SR2B_2/dff3B_0/D SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Smb SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M1375 SubB_0/SR2B_2/dff3B_0/D SS0 SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M1376 SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Min1 nor2_0/out SubB_0/abs_0/sum Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=85p ps=54u 
M1377 SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Min1 SubB_0/SR2B_2/mux4x1_0/mux2x1_1/Smb SubB_0/abs_0/sum Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1378 SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Min1 SubB_0/SR2B_2/mux4x1_0/mux2x1_1/Smb D0 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M1379 SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Min1 nor2_0/out D0 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M1380 SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Smb SS0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1381 SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Smb SS0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1382 SubB_0/SR2B_2/mux4x1_0/mux2x1_1/Smb nor2_0/out Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1383 SubB_0/SR2B_2/mux4x1_0/mux2x1_1/Smb nor2_0/out GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1384 SubB_0/SR2B_1/dff3B_7/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1385 SubB_0/SR2B_1/dff3B_7/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1386 SubB_0/SR2B_1/dff3B_7/gate_0/S SubB_0/SR2B_1/dff3B_7/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1387 SubB_0/SR2B_1/dff3B_7/gate_0/S SubB_0/SR2B_1/dff3B_7/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1388 SubB_0/SR2B_1/dff3B_7/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1389 SubB_0/SR2B_1/dff3B_7/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1390 SubB_0/SR2B_1/dff3B_7/gate_3/Gout SubB_0/SR2B_1/Q7 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1391 SubB_0/SR2B_1/dff3B_7/gate_3/Gout SubB_0/SR2B_1/Q7 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1392 SubB_0/SR2B_1/dff3B_7/gate_3/Gout fsm_0/CLK SubB_0/SR2B_1/dff3B_7/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1393 SubB_0/SR2B_1/dff3B_7/gate_3/Gout SubB_0/SR2B_1/dff3B_7/gate_1/S SubB_0/SR2B_1/dff3B_7/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1394 SubB_0/SR2B_1/dff3B_7/gate_2/Gout SubB_0/SR2B_1/dff3B_7/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1395 SubB_0/SR2B_1/dff3B_7/gate_2/Gout SubB_0/SR2B_1/dff3B_7/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1396 SubB_0/SR2B_1/dff3B_7/gate_2/Gout SubB_0/SR2B_1/dff3B_7/gate_2/S SubB_0/SR2B_1/dff3B_7/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1397 SubB_0/SR2B_1/dff3B_7/gate_2/Gout SubB_0/SR2B_1/dff3B_7/gate_0/S SubB_0/SR2B_1/dff3B_7/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1398 SubB_0/SR2B_1/dff3B_7/Qb SubB_0/SR2B_1/Q7 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1399 SubB_0/SR2B_1/dff3B_7/Qb SubB_0/SR2B_1/Q7 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1400 SubB_0/SR2B_1/Q7 SubB_0/SR2B_1/dff3B_7/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=124p pd=82u as=0p ps=0u 
M1401 SubB_0/SR2B_1/Q7 SubB_0/SR2B_1/dff3B_7/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=75p pd=66u as=0p ps=0u 
M1402 SubB_0/SR2B_1/dff3B_7/gate_3/Gin SubB_0/SR2B_1/dff3B_7/gate_1/S SubB_0/SR2B_1/dff3B_7/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1403 SubB_0/SR2B_1/dff3B_7/gate_3/Gin fsm_0/CLK SubB_0/SR2B_1/dff3B_7/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1404 SubB_0/SR2B_1/dff3B_7/gate_1/Gin SubB_0/SR2B_1/dff3B_7/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1405 SubB_0/SR2B_1/dff3B_7/gate_1/Gin SubB_0/SR2B_1/dff3B_7/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1406 SubB_0/SR2B_1/dff3B_7/gate_2/Gin SubB_0/SR2B_1/dff3B_7/gate_0/S SubB_0/SR2B_1/dff3B_7/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1407 SubB_0/SR2B_1/dff3B_7/gate_2/Gin SubB_0/SR2B_1/dff3B_7/gate_2/S SubB_0/SR2B_1/dff3B_7/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1408 SubB_0/SR2B_1/dff3B_7/gate_0/Gin SubB_0/SR2B_1/dff3B_7/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1409 SubB_0/SR2B_1/dff3B_7/gate_0/Gin SubB_0/SR2B_1/dff3B_7/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1410 SubB_0/SR2B_1/dff3B_7/inverter_11/in SubB_0/SR2B_1/dff3B_7/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1411 Vdd SubB_0/SR2B_1/dff3B_7/D SubB_0/SR2B_1/dff3B_7/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1412 SubB_0/SR2B_1/dff3B_7/nand2_0/a_n37_n6# SubB_0/SR2B_1/dff3B_7/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1413 SubB_0/SR2B_1/dff3B_7/inverter_11/in SubB_0/SR2B_1/dff3B_7/D SubB_0/SR2B_1/dff3B_7/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1414 SubB_0/SR2B_1/dff3B_7/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1415 SubB_0/SR2B_1/dff3B_7/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1416 SubB_0/SR2B_1/dff3B_6/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1417 SubB_0/SR2B_1/dff3B_6/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1418 SubB_0/SR2B_1/dff3B_6/gate_0/S SubB_0/SR2B_1/dff3B_6/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1419 SubB_0/SR2B_1/dff3B_6/gate_0/S SubB_0/SR2B_1/dff3B_6/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1420 SubB_0/SR2B_1/dff3B_6/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1421 SubB_0/SR2B_1/dff3B_6/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1422 SubB_0/SR2B_1/dff3B_6/gate_3/Gout SubB_0/SR2B_1/Q6 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1423 SubB_0/SR2B_1/dff3B_6/gate_3/Gout SubB_0/SR2B_1/Q6 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1424 SubB_0/SR2B_1/dff3B_6/gate_3/Gout fsm_0/CLK SubB_0/SR2B_1/dff3B_6/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1425 SubB_0/SR2B_1/dff3B_6/gate_3/Gout SubB_0/SR2B_1/dff3B_6/gate_1/S SubB_0/SR2B_1/dff3B_6/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1426 SubB_0/SR2B_1/dff3B_6/gate_2/Gout SubB_0/SR2B_1/dff3B_6/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1427 SubB_0/SR2B_1/dff3B_6/gate_2/Gout SubB_0/SR2B_1/dff3B_6/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1428 SubB_0/SR2B_1/dff3B_6/gate_2/Gout SubB_0/SR2B_1/dff3B_6/gate_2/S SubB_0/SR2B_1/dff3B_6/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1429 SubB_0/SR2B_1/dff3B_6/gate_2/Gout SubB_0/SR2B_1/dff3B_6/gate_0/S SubB_0/SR2B_1/dff3B_6/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1430 SubB_0/SR2B_1/dff3B_6/Qb SubB_0/SR2B_1/Q6 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1431 SubB_0/SR2B_1/dff3B_6/Qb SubB_0/SR2B_1/Q6 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1432 SubB_0/SR2B_1/Q6 SubB_0/SR2B_1/dff3B_6/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M1433 SubB_0/SR2B_1/Q6 SubB_0/SR2B_1/dff3B_6/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M1434 SubB_0/SR2B_1/dff3B_6/gate_3/Gin SubB_0/SR2B_1/dff3B_6/gate_1/S SubB_0/SR2B_1/dff3B_6/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1435 SubB_0/SR2B_1/dff3B_6/gate_3/Gin fsm_0/CLK SubB_0/SR2B_1/dff3B_6/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1436 SubB_0/SR2B_1/dff3B_6/gate_1/Gin SubB_0/SR2B_1/dff3B_6/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1437 SubB_0/SR2B_1/dff3B_6/gate_1/Gin SubB_0/SR2B_1/dff3B_6/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1438 SubB_0/SR2B_1/dff3B_6/gate_2/Gin SubB_0/SR2B_1/dff3B_6/gate_0/S SubB_0/SR2B_1/dff3B_6/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1439 SubB_0/SR2B_1/dff3B_6/gate_2/Gin SubB_0/SR2B_1/dff3B_6/gate_2/S SubB_0/SR2B_1/dff3B_6/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1440 SubB_0/SR2B_1/dff3B_6/gate_0/Gin SubB_0/SR2B_1/dff3B_6/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1441 SubB_0/SR2B_1/dff3B_6/gate_0/Gin SubB_0/SR2B_1/dff3B_6/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1442 SubB_0/SR2B_1/dff3B_6/inverter_11/in SubB_0/SR2B_1/dff3B_6/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1443 Vdd SubB_0/SR2B_1/dff3B_6/D SubB_0/SR2B_1/dff3B_6/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1444 SubB_0/SR2B_1/dff3B_6/nand2_0/a_n37_n6# SubB_0/SR2B_1/dff3B_6/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1445 SubB_0/SR2B_1/dff3B_6/inverter_11/in SubB_0/SR2B_1/dff3B_6/D SubB_0/SR2B_1/dff3B_6/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1446 SubB_0/SR2B_1/dff3B_6/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1447 SubB_0/SR2B_1/dff3B_6/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1448 SubB_0/SR2B_1/dff3B_5/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1449 SubB_0/SR2B_1/dff3B_5/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1450 SubB_0/SR2B_1/dff3B_5/gate_0/S SubB_0/SR2B_1/dff3B_5/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1451 SubB_0/SR2B_1/dff3B_5/gate_0/S SubB_0/SR2B_1/dff3B_5/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1452 SubB_0/SR2B_1/dff3B_5/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1453 SubB_0/SR2B_1/dff3B_5/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1454 SubB_0/SR2B_1/dff3B_5/gate_3/Gout SubB_0/SR2B_1/Q5 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1455 SubB_0/SR2B_1/dff3B_5/gate_3/Gout SubB_0/SR2B_1/Q5 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1456 SubB_0/SR2B_1/dff3B_5/gate_3/Gout fsm_0/CLK SubB_0/SR2B_1/dff3B_5/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1457 SubB_0/SR2B_1/dff3B_5/gate_3/Gout SubB_0/SR2B_1/dff3B_5/gate_1/S SubB_0/SR2B_1/dff3B_5/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1458 SubB_0/SR2B_1/dff3B_5/gate_2/Gout SubB_0/SR2B_1/dff3B_5/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1459 SubB_0/SR2B_1/dff3B_5/gate_2/Gout SubB_0/SR2B_1/dff3B_5/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1460 SubB_0/SR2B_1/dff3B_5/gate_2/Gout SubB_0/SR2B_1/dff3B_5/gate_2/S SubB_0/SR2B_1/dff3B_5/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1461 SubB_0/SR2B_1/dff3B_5/gate_2/Gout SubB_0/SR2B_1/dff3B_5/gate_0/S SubB_0/SR2B_1/dff3B_5/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1462 SubB_0/SR2B_1/dff3B_5/Qb SubB_0/SR2B_1/Q5 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1463 SubB_0/SR2B_1/dff3B_5/Qb SubB_0/SR2B_1/Q5 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1464 SubB_0/SR2B_1/Q5 SubB_0/SR2B_1/dff3B_5/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M1465 SubB_0/SR2B_1/Q5 SubB_0/SR2B_1/dff3B_5/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M1466 SubB_0/SR2B_1/dff3B_5/gate_3/Gin SubB_0/SR2B_1/dff3B_5/gate_1/S SubB_0/SR2B_1/dff3B_5/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1467 SubB_0/SR2B_1/dff3B_5/gate_3/Gin fsm_0/CLK SubB_0/SR2B_1/dff3B_5/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1468 SubB_0/SR2B_1/dff3B_5/gate_1/Gin SubB_0/SR2B_1/dff3B_5/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1469 SubB_0/SR2B_1/dff3B_5/gate_1/Gin SubB_0/SR2B_1/dff3B_5/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1470 SubB_0/SR2B_1/dff3B_5/gate_2/Gin SubB_0/SR2B_1/dff3B_5/gate_0/S SubB_0/SR2B_1/dff3B_5/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1471 SubB_0/SR2B_1/dff3B_5/gate_2/Gin SubB_0/SR2B_1/dff3B_5/gate_2/S SubB_0/SR2B_1/dff3B_5/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1472 SubB_0/SR2B_1/dff3B_5/gate_0/Gin SubB_0/SR2B_1/dff3B_5/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1473 SubB_0/SR2B_1/dff3B_5/gate_0/Gin SubB_0/SR2B_1/dff3B_5/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1474 SubB_0/SR2B_1/dff3B_5/inverter_11/in SubB_0/SR2B_1/dff3B_5/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1475 Vdd SubB_0/SR2B_1/dff3B_5/D SubB_0/SR2B_1/dff3B_5/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1476 SubB_0/SR2B_1/dff3B_5/nand2_0/a_n37_n6# SubB_0/SR2B_1/dff3B_5/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1477 SubB_0/SR2B_1/dff3B_5/inverter_11/in SubB_0/SR2B_1/dff3B_5/D SubB_0/SR2B_1/dff3B_5/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1478 SubB_0/SR2B_1/dff3B_5/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1479 SubB_0/SR2B_1/dff3B_5/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1480 SubB_0/SR2B_1/dff3B_4/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1481 SubB_0/SR2B_1/dff3B_4/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1482 SubB_0/SR2B_1/dff3B_4/gate_0/S SubB_0/SR2B_1/dff3B_4/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1483 SubB_0/SR2B_1/dff3B_4/gate_0/S SubB_0/SR2B_1/dff3B_4/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1484 SubB_0/SR2B_1/dff3B_4/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1485 SubB_0/SR2B_1/dff3B_4/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1486 SubB_0/SR2B_1/dff3B_4/gate_3/Gout SubB_0/SR2B_1/Q4 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1487 SubB_0/SR2B_1/dff3B_4/gate_3/Gout SubB_0/SR2B_1/Q4 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1488 SubB_0/SR2B_1/dff3B_4/gate_3/Gout fsm_0/CLK SubB_0/SR2B_1/dff3B_4/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1489 SubB_0/SR2B_1/dff3B_4/gate_3/Gout SubB_0/SR2B_1/dff3B_4/gate_1/S SubB_0/SR2B_1/dff3B_4/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1490 SubB_0/SR2B_1/dff3B_4/gate_2/Gout SubB_0/SR2B_1/dff3B_4/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1491 SubB_0/SR2B_1/dff3B_4/gate_2/Gout SubB_0/SR2B_1/dff3B_4/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1492 SubB_0/SR2B_1/dff3B_4/gate_2/Gout SubB_0/SR2B_1/dff3B_4/gate_2/S SubB_0/SR2B_1/dff3B_4/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1493 SubB_0/SR2B_1/dff3B_4/gate_2/Gout SubB_0/SR2B_1/dff3B_4/gate_0/S SubB_0/SR2B_1/dff3B_4/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1494 SubB_0/SR2B_1/dff3B_4/Qb SubB_0/SR2B_1/Q4 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1495 SubB_0/SR2B_1/dff3B_4/Qb SubB_0/SR2B_1/Q4 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1496 SubB_0/SR2B_1/Q4 SubB_0/SR2B_1/dff3B_4/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M1497 SubB_0/SR2B_1/Q4 SubB_0/SR2B_1/dff3B_4/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M1498 SubB_0/SR2B_1/dff3B_4/gate_3/Gin SubB_0/SR2B_1/dff3B_4/gate_1/S SubB_0/SR2B_1/dff3B_4/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1499 SubB_0/SR2B_1/dff3B_4/gate_3/Gin fsm_0/CLK SubB_0/SR2B_1/dff3B_4/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1500 SubB_0/SR2B_1/dff3B_4/gate_1/Gin SubB_0/SR2B_1/dff3B_4/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1501 SubB_0/SR2B_1/dff3B_4/gate_1/Gin SubB_0/SR2B_1/dff3B_4/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1502 SubB_0/SR2B_1/dff3B_4/gate_2/Gin SubB_0/SR2B_1/dff3B_4/gate_0/S SubB_0/SR2B_1/dff3B_4/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1503 SubB_0/SR2B_1/dff3B_4/gate_2/Gin SubB_0/SR2B_1/dff3B_4/gate_2/S SubB_0/SR2B_1/dff3B_4/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1504 SubB_0/SR2B_1/dff3B_4/gate_0/Gin SubB_0/SR2B_1/dff3B_4/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1505 SubB_0/SR2B_1/dff3B_4/gate_0/Gin SubB_0/SR2B_1/dff3B_4/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1506 SubB_0/SR2B_1/dff3B_4/inverter_11/in SubB_0/SR2B_1/dff3B_4/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1507 Vdd SubB_0/SR2B_1/dff3B_4/D SubB_0/SR2B_1/dff3B_4/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1508 SubB_0/SR2B_1/dff3B_4/nand2_0/a_n37_n6# SubB_0/SR2B_1/dff3B_4/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1509 SubB_0/SR2B_1/dff3B_4/inverter_11/in SubB_0/SR2B_1/dff3B_4/D SubB_0/SR2B_1/dff3B_4/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1510 SubB_0/SR2B_1/dff3B_4/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1511 SubB_0/SR2B_1/dff3B_4/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1512 SubB_0/SR2B_1/dff3B_3/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1513 SubB_0/SR2B_1/dff3B_3/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1514 SubB_0/SR2B_1/dff3B_3/gate_0/S SubB_0/SR2B_1/dff3B_3/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1515 SubB_0/SR2B_1/dff3B_3/gate_0/S SubB_0/SR2B_1/dff3B_3/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1516 SubB_0/SR2B_1/dff3B_3/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1517 SubB_0/SR2B_1/dff3B_3/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1518 SubB_0/SR2B_1/dff3B_3/gate_3/Gout SubB_0/SR2B_1/Q3 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1519 SubB_0/SR2B_1/dff3B_3/gate_3/Gout SubB_0/SR2B_1/Q3 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1520 SubB_0/SR2B_1/dff3B_3/gate_3/Gout fsm_0/CLK SubB_0/SR2B_1/dff3B_3/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1521 SubB_0/SR2B_1/dff3B_3/gate_3/Gout SubB_0/SR2B_1/dff3B_3/gate_1/S SubB_0/SR2B_1/dff3B_3/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1522 SubB_0/SR2B_1/dff3B_3/gate_2/Gout SubB_0/SR2B_1/dff3B_3/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1523 SubB_0/SR2B_1/dff3B_3/gate_2/Gout SubB_0/SR2B_1/dff3B_3/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1524 SubB_0/SR2B_1/dff3B_3/gate_2/Gout SubB_0/SR2B_1/dff3B_3/gate_2/S SubB_0/SR2B_1/dff3B_3/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1525 SubB_0/SR2B_1/dff3B_3/gate_2/Gout SubB_0/SR2B_1/dff3B_3/gate_0/S SubB_0/SR2B_1/dff3B_3/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1526 SubB_0/SR2B_1/dff3B_3/Qb SubB_0/SR2B_1/Q3 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1527 SubB_0/SR2B_1/dff3B_3/Qb SubB_0/SR2B_1/Q3 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1528 SubB_0/SR2B_1/Q3 SubB_0/SR2B_1/dff3B_3/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M1529 SubB_0/SR2B_1/Q3 SubB_0/SR2B_1/dff3B_3/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M1530 SubB_0/SR2B_1/dff3B_3/gate_3/Gin SubB_0/SR2B_1/dff3B_3/gate_1/S SubB_0/SR2B_1/dff3B_3/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1531 SubB_0/SR2B_1/dff3B_3/gate_3/Gin fsm_0/CLK SubB_0/SR2B_1/dff3B_3/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1532 SubB_0/SR2B_1/dff3B_3/gate_1/Gin SubB_0/SR2B_1/dff3B_3/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1533 SubB_0/SR2B_1/dff3B_3/gate_1/Gin SubB_0/SR2B_1/dff3B_3/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1534 SubB_0/SR2B_1/dff3B_3/gate_2/Gin SubB_0/SR2B_1/dff3B_3/gate_0/S SubB_0/SR2B_1/dff3B_3/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1535 SubB_0/SR2B_1/dff3B_3/gate_2/Gin SubB_0/SR2B_1/dff3B_3/gate_2/S SubB_0/SR2B_1/dff3B_3/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1536 SubB_0/SR2B_1/dff3B_3/gate_0/Gin SubB_0/SR2B_1/dff3B_3/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1537 SubB_0/SR2B_1/dff3B_3/gate_0/Gin SubB_0/SR2B_1/dff3B_3/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1538 SubB_0/SR2B_1/dff3B_3/inverter_11/in SubB_0/SR2B_1/dff3B_3/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1539 Vdd SubB_0/SR2B_1/dff3B_3/D SubB_0/SR2B_1/dff3B_3/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1540 SubB_0/SR2B_1/dff3B_3/nand2_0/a_n37_n6# SubB_0/SR2B_1/dff3B_3/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1541 SubB_0/SR2B_1/dff3B_3/inverter_11/in SubB_0/SR2B_1/dff3B_3/D SubB_0/SR2B_1/dff3B_3/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1542 SubB_0/SR2B_1/dff3B_3/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1543 SubB_0/SR2B_1/dff3B_3/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1544 SubB_0/SR2B_1/dff3B_2/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1545 SubB_0/SR2B_1/dff3B_2/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1546 SubB_0/SR2B_1/dff3B_2/gate_0/S SubB_0/SR2B_1/dff3B_2/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1547 SubB_0/SR2B_1/dff3B_2/gate_0/S SubB_0/SR2B_1/dff3B_2/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1548 SubB_0/SR2B_1/dff3B_2/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1549 SubB_0/SR2B_1/dff3B_2/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1550 SubB_0/SR2B_1/dff3B_2/gate_3/Gout SubB_0/SR2B_1/Q2 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1551 SubB_0/SR2B_1/dff3B_2/gate_3/Gout SubB_0/SR2B_1/Q2 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1552 SubB_0/SR2B_1/dff3B_2/gate_3/Gout fsm_0/CLK SubB_0/SR2B_1/dff3B_2/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1553 SubB_0/SR2B_1/dff3B_2/gate_3/Gout SubB_0/SR2B_1/dff3B_2/gate_1/S SubB_0/SR2B_1/dff3B_2/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1554 SubB_0/SR2B_1/dff3B_2/gate_2/Gout SubB_0/SR2B_1/dff3B_2/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1555 SubB_0/SR2B_1/dff3B_2/gate_2/Gout SubB_0/SR2B_1/dff3B_2/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1556 SubB_0/SR2B_1/dff3B_2/gate_2/Gout SubB_0/SR2B_1/dff3B_2/gate_2/S SubB_0/SR2B_1/dff3B_2/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1557 SubB_0/SR2B_1/dff3B_2/gate_2/Gout SubB_0/SR2B_1/dff3B_2/gate_0/S SubB_0/SR2B_1/dff3B_2/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1558 SubB_0/SR2B_1/dff3B_2/Qb SubB_0/SR2B_1/Q2 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1559 SubB_0/SR2B_1/dff3B_2/Qb SubB_0/SR2B_1/Q2 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1560 SubB_0/SR2B_1/Q2 SubB_0/SR2B_1/dff3B_2/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M1561 SubB_0/SR2B_1/Q2 SubB_0/SR2B_1/dff3B_2/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M1562 SubB_0/SR2B_1/dff3B_2/gate_3/Gin SubB_0/SR2B_1/dff3B_2/gate_1/S SubB_0/SR2B_1/dff3B_2/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1563 SubB_0/SR2B_1/dff3B_2/gate_3/Gin fsm_0/CLK SubB_0/SR2B_1/dff3B_2/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1564 SubB_0/SR2B_1/dff3B_2/gate_1/Gin SubB_0/SR2B_1/dff3B_2/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1565 SubB_0/SR2B_1/dff3B_2/gate_1/Gin SubB_0/SR2B_1/dff3B_2/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1566 SubB_0/SR2B_1/dff3B_2/gate_2/Gin SubB_0/SR2B_1/dff3B_2/gate_0/S SubB_0/SR2B_1/dff3B_2/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1567 SubB_0/SR2B_1/dff3B_2/gate_2/Gin SubB_0/SR2B_1/dff3B_2/gate_2/S SubB_0/SR2B_1/dff3B_2/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1568 SubB_0/SR2B_1/dff3B_2/gate_0/Gin SubB_0/SR2B_1/dff3B_2/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1569 SubB_0/SR2B_1/dff3B_2/gate_0/Gin SubB_0/SR2B_1/dff3B_2/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1570 SubB_0/SR2B_1/dff3B_2/inverter_11/in SubB_0/SR2B_1/dff3B_2/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1571 Vdd SubB_0/SR2B_1/dff3B_2/D SubB_0/SR2B_1/dff3B_2/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1572 SubB_0/SR2B_1/dff3B_2/nand2_0/a_n37_n6# SubB_0/SR2B_1/dff3B_2/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1573 SubB_0/SR2B_1/dff3B_2/inverter_11/in SubB_0/SR2B_1/dff3B_2/D SubB_0/SR2B_1/dff3B_2/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1574 SubB_0/SR2B_1/dff3B_2/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1575 SubB_0/SR2B_1/dff3B_2/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1576 SubB_0/SR2B_1/dff3B_1/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1577 SubB_0/SR2B_1/dff3B_1/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1578 SubB_0/SR2B_1/dff3B_1/gate_0/S SubB_0/SR2B_1/dff3B_1/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1579 SubB_0/SR2B_1/dff3B_1/gate_0/S SubB_0/SR2B_1/dff3B_1/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1580 SubB_0/SR2B_1/dff3B_1/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1581 SubB_0/SR2B_1/dff3B_1/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1582 SubB_0/SR2B_1/dff3B_1/gate_3/Gout SubB_0/SR2B_1/Q1 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1583 SubB_0/SR2B_1/dff3B_1/gate_3/Gout SubB_0/SR2B_1/Q1 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1584 SubB_0/SR2B_1/dff3B_1/gate_3/Gout fsm_0/CLK SubB_0/SR2B_1/dff3B_1/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1585 SubB_0/SR2B_1/dff3B_1/gate_3/Gout SubB_0/SR2B_1/dff3B_1/gate_1/S SubB_0/SR2B_1/dff3B_1/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1586 SubB_0/SR2B_1/dff3B_1/gate_2/Gout SubB_0/SR2B_1/dff3B_1/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1587 SubB_0/SR2B_1/dff3B_1/gate_2/Gout SubB_0/SR2B_1/dff3B_1/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1588 SubB_0/SR2B_1/dff3B_1/gate_2/Gout SubB_0/SR2B_1/dff3B_1/gate_2/S SubB_0/SR2B_1/dff3B_1/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1589 SubB_0/SR2B_1/dff3B_1/gate_2/Gout SubB_0/SR2B_1/dff3B_1/gate_0/S SubB_0/SR2B_1/dff3B_1/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1590 SubB_0/SR2B_1/dff3B_1/Qb SubB_0/SR2B_1/Q1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1591 SubB_0/SR2B_1/dff3B_1/Qb SubB_0/SR2B_1/Q1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1592 SubB_0/SR2B_1/Q1 SubB_0/SR2B_1/dff3B_1/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M1593 SubB_0/SR2B_1/Q1 SubB_0/SR2B_1/dff3B_1/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M1594 SubB_0/SR2B_1/dff3B_1/gate_3/Gin SubB_0/SR2B_1/dff3B_1/gate_1/S SubB_0/SR2B_1/dff3B_1/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1595 SubB_0/SR2B_1/dff3B_1/gate_3/Gin fsm_0/CLK SubB_0/SR2B_1/dff3B_1/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1596 SubB_0/SR2B_1/dff3B_1/gate_1/Gin SubB_0/SR2B_1/dff3B_1/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1597 SubB_0/SR2B_1/dff3B_1/gate_1/Gin SubB_0/SR2B_1/dff3B_1/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1598 SubB_0/SR2B_1/dff3B_1/gate_2/Gin SubB_0/SR2B_1/dff3B_1/gate_0/S SubB_0/SR2B_1/dff3B_1/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1599 SubB_0/SR2B_1/dff3B_1/gate_2/Gin SubB_0/SR2B_1/dff3B_1/gate_2/S SubB_0/SR2B_1/dff3B_1/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1600 SubB_0/SR2B_1/dff3B_1/gate_0/Gin SubB_0/SR2B_1/dff3B_1/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1601 SubB_0/SR2B_1/dff3B_1/gate_0/Gin SubB_0/SR2B_1/dff3B_1/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1602 SubB_0/SR2B_1/dff3B_1/inverter_11/in SubB_0/SR2B_1/dff3B_1/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1603 Vdd SubB_0/SR2B_1/dff3B_1/D SubB_0/SR2B_1/dff3B_1/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1604 SubB_0/SR2B_1/dff3B_1/nand2_0/a_n37_n6# SubB_0/SR2B_1/dff3B_1/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1605 SubB_0/SR2B_1/dff3B_1/inverter_11/in SubB_0/SR2B_1/dff3B_1/D SubB_0/SR2B_1/dff3B_1/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1606 SubB_0/SR2B_1/dff3B_1/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1607 SubB_0/SR2B_1/dff3B_1/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1608 SubB_0/SR2B_1/dff3B_0/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1609 SubB_0/SR2B_1/dff3B_0/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1610 SubB_0/SR2B_1/dff3B_0/gate_0/S SubB_0/SR2B_1/dff3B_0/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1611 SubB_0/SR2B_1/dff3B_0/gate_0/S SubB_0/SR2B_1/dff3B_0/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1612 SubB_0/SR2B_1/dff3B_0/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1613 SubB_0/SR2B_1/dff3B_0/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1614 SubB_0/SR2B_1/dff3B_0/gate_3/Gout SubB_0/QB0 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1615 SubB_0/SR2B_1/dff3B_0/gate_3/Gout SubB_0/QB0 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1616 SubB_0/SR2B_1/dff3B_0/gate_3/Gout fsm_0/CLK SubB_0/SR2B_1/dff3B_0/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1617 SubB_0/SR2B_1/dff3B_0/gate_3/Gout SubB_0/SR2B_1/dff3B_0/gate_1/S SubB_0/SR2B_1/dff3B_0/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1618 SubB_0/SR2B_1/dff3B_0/gate_2/Gout SubB_0/SR2B_1/dff3B_0/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1619 SubB_0/SR2B_1/dff3B_0/gate_2/Gout SubB_0/SR2B_1/dff3B_0/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1620 SubB_0/SR2B_1/dff3B_0/gate_2/Gout SubB_0/SR2B_1/dff3B_0/gate_2/S SubB_0/SR2B_1/dff3B_0/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1621 SubB_0/SR2B_1/dff3B_0/gate_2/Gout SubB_0/SR2B_1/dff3B_0/gate_0/S SubB_0/SR2B_1/dff3B_0/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1622 SubB_0/SR2B_1/dff3B_0/Qb SubB_0/QB0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1623 SubB_0/SR2B_1/dff3B_0/Qb SubB_0/QB0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1624 SubB_0/QB0 SubB_0/SR2B_1/dff3B_0/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M1625 SubB_0/QB0 SubB_0/SR2B_1/dff3B_0/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M1626 SubB_0/SR2B_1/dff3B_0/gate_3/Gin SubB_0/SR2B_1/dff3B_0/gate_1/S SubB_0/SR2B_1/dff3B_0/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1627 SubB_0/SR2B_1/dff3B_0/gate_3/Gin fsm_0/CLK SubB_0/SR2B_1/dff3B_0/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1628 SubB_0/SR2B_1/dff3B_0/gate_1/Gin SubB_0/SR2B_1/dff3B_0/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1629 SubB_0/SR2B_1/dff3B_0/gate_1/Gin SubB_0/SR2B_1/dff3B_0/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1630 SubB_0/SR2B_1/dff3B_0/gate_2/Gin SubB_0/SR2B_1/dff3B_0/gate_0/S SubB_0/SR2B_1/dff3B_0/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1631 SubB_0/SR2B_1/dff3B_0/gate_2/Gin SubB_0/SR2B_1/dff3B_0/gate_2/S SubB_0/SR2B_1/dff3B_0/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1632 SubB_0/SR2B_1/dff3B_0/gate_0/Gin SubB_0/SR2B_1/dff3B_0/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1633 SubB_0/SR2B_1/dff3B_0/gate_0/Gin SubB_0/SR2B_1/dff3B_0/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1634 SubB_0/SR2B_1/dff3B_0/inverter_11/in SubB_0/SR2B_1/dff3B_0/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1635 Vdd SubB_0/SR2B_1/dff3B_0/D SubB_0/SR2B_1/dff3B_0/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1636 SubB_0/SR2B_1/dff3B_0/nand2_0/a_n37_n6# SubB_0/SR2B_1/dff3B_0/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1637 SubB_0/SR2B_1/dff3B_0/inverter_11/in SubB_0/SR2B_1/dff3B_0/D SubB_0/SR2B_1/dff3B_0/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1638 SubB_0/SR2B_1/dff3B_0/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1639 SubB_0/SR2B_1/dff3B_0/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1640 SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Min2 SB1 SubB_0/SR2B_1/Q7 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M1641 SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Min2 SubB_0/SR2B_1/mux4x1_7/mux2x1_1/Smb SubB_0/SR2B_1/Q7 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M1642 SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Min2 SubB_0/SR2B_1/mux4x1_7/mux2x1_1/Smb SubB_0/QB0 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1643 SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Min2 SB1 SubB_0/QB0 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1644 SubB_0/SR2B_1/dff3B_7/D SB0 SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M1645 SubB_0/SR2B_1/dff3B_7/D SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Smb SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M1646 SubB_0/SR2B_1/dff3B_7/D SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Smb SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M1647 SubB_0/SR2B_1/dff3B_7/D SB0 SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M1648 SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Min1 SB1 SubB_0/SR2B_1/Q6 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1649 SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Min1 SubB_0/SR2B_1/mux4x1_7/mux2x1_1/Smb SubB_0/SR2B_1/Q6 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1650 SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Min1 SubB_0/SR2B_1/mux4x1_7/mux2x1_1/Smb B7 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M1651 SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Min1 SB1 B7 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M1652 SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Smb SB0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1653 SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Smb SB0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1654 SubB_0/SR2B_1/mux4x1_7/mux2x1_1/Smb SB1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1655 SubB_0/SR2B_1/mux4x1_7/mux2x1_1/Smb SB1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1656 SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Min2 SB1 SubB_0/SR2B_1/Q6 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M1657 SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Min2 SubB_0/SR2B_1/mux4x1_6/mux2x1_1/Smb SubB_0/SR2B_1/Q6 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M1658 SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Min2 SubB_0/SR2B_1/mux4x1_6/mux2x1_1/Smb SubB_0/SR2B_1/Q7 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1659 SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Min2 SB1 SubB_0/SR2B_1/Q7 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1660 SubB_0/SR2B_1/dff3B_6/D SB0 SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M1661 SubB_0/SR2B_1/dff3B_6/D SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Smb SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M1662 SubB_0/SR2B_1/dff3B_6/D SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Smb SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M1663 SubB_0/SR2B_1/dff3B_6/D SB0 SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M1664 SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Min1 SB1 SubB_0/SR2B_1/Q5 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1665 SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Min1 SubB_0/SR2B_1/mux4x1_6/mux2x1_1/Smb SubB_0/SR2B_1/Q5 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1666 SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Min1 SubB_0/SR2B_1/mux4x1_6/mux2x1_1/Smb B6 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M1667 SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Min1 SB1 B6 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M1668 SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Smb SB0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1669 SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Smb SB0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1670 SubB_0/SR2B_1/mux4x1_6/mux2x1_1/Smb SB1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1671 SubB_0/SR2B_1/mux4x1_6/mux2x1_1/Smb SB1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1672 SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Min2 SB1 SubB_0/SR2B_1/Q5 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M1673 SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Min2 SubB_0/SR2B_1/mux4x1_5/mux2x1_1/Smb SubB_0/SR2B_1/Q5 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M1674 SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Min2 SubB_0/SR2B_1/mux4x1_5/mux2x1_1/Smb SubB_0/SR2B_1/Q6 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1675 SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Min2 SB1 SubB_0/SR2B_1/Q6 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1676 SubB_0/SR2B_1/dff3B_5/D SB0 SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M1677 SubB_0/SR2B_1/dff3B_5/D SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Smb SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M1678 SubB_0/SR2B_1/dff3B_5/D SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Smb SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M1679 SubB_0/SR2B_1/dff3B_5/D SB0 SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M1680 SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Min1 SB1 SubB_0/SR2B_1/Q4 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1681 SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Min1 SubB_0/SR2B_1/mux4x1_5/mux2x1_1/Smb SubB_0/SR2B_1/Q4 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1682 SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Min1 SubB_0/SR2B_1/mux4x1_5/mux2x1_1/Smb B5 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M1683 SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Min1 SB1 B5 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M1684 SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Smb SB0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1685 SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Smb SB0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1686 SubB_0/SR2B_1/mux4x1_5/mux2x1_1/Smb SB1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1687 SubB_0/SR2B_1/mux4x1_5/mux2x1_1/Smb SB1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1688 SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Min2 SB1 SubB_0/SR2B_1/Q4 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M1689 SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Min2 SubB_0/SR2B_1/mux4x1_4/mux2x1_1/Smb SubB_0/SR2B_1/Q4 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M1690 SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Min2 SubB_0/SR2B_1/mux4x1_4/mux2x1_1/Smb SubB_0/SR2B_1/Q5 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1691 SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Min2 SB1 SubB_0/SR2B_1/Q5 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1692 SubB_0/SR2B_1/dff3B_4/D SB0 SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M1693 SubB_0/SR2B_1/dff3B_4/D SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Smb SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M1694 SubB_0/SR2B_1/dff3B_4/D SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Smb SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M1695 SubB_0/SR2B_1/dff3B_4/D SB0 SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M1696 SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Min1 SB1 SubB_0/SR2B_1/Q3 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1697 SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Min1 SubB_0/SR2B_1/mux4x1_4/mux2x1_1/Smb SubB_0/SR2B_1/Q3 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1698 SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Min1 SubB_0/SR2B_1/mux4x1_4/mux2x1_1/Smb B4 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M1699 SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Min1 SB1 B4 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M1700 SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Smb SB0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1701 SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Smb SB0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1702 SubB_0/SR2B_1/mux4x1_4/mux2x1_1/Smb SB1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1703 SubB_0/SR2B_1/mux4x1_4/mux2x1_1/Smb SB1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1704 SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Min2 SB1 SubB_0/SR2B_1/Q3 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M1705 SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Min2 SubB_0/SR2B_1/mux4x1_3/mux2x1_1/Smb SubB_0/SR2B_1/Q3 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M1706 SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Min2 SubB_0/SR2B_1/mux4x1_3/mux2x1_1/Smb SubB_0/SR2B_1/Q4 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1707 SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Min2 SB1 SubB_0/SR2B_1/Q4 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1708 SubB_0/SR2B_1/dff3B_3/D SB0 SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M1709 SubB_0/SR2B_1/dff3B_3/D SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Smb SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M1710 SubB_0/SR2B_1/dff3B_3/D SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Smb SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M1711 SubB_0/SR2B_1/dff3B_3/D SB0 SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M1712 SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Min1 SB1 SubB_0/SR2B_1/Q2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1713 SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Min1 SubB_0/SR2B_1/mux4x1_3/mux2x1_1/Smb SubB_0/SR2B_1/Q2 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1714 SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Min1 SubB_0/SR2B_1/mux4x1_3/mux2x1_1/Smb B3 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M1715 SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Min1 SB1 B3 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M1716 SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Smb SB0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1717 SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Smb SB0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1718 SubB_0/SR2B_1/mux4x1_3/mux2x1_1/Smb SB1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1719 SubB_0/SR2B_1/mux4x1_3/mux2x1_1/Smb SB1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1720 SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Min2 SB1 SubB_0/SR2B_1/Q2 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M1721 SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Min2 SubB_0/SR2B_1/mux4x1_2/mux2x1_1/Smb SubB_0/SR2B_1/Q2 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M1722 SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Min2 SubB_0/SR2B_1/mux4x1_2/mux2x1_1/Smb SubB_0/SR2B_1/Q3 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1723 SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Min2 SB1 SubB_0/SR2B_1/Q3 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1724 SubB_0/SR2B_1/dff3B_2/D SB0 SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M1725 SubB_0/SR2B_1/dff3B_2/D SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Smb SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M1726 SubB_0/SR2B_1/dff3B_2/D SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Smb SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M1727 SubB_0/SR2B_1/dff3B_2/D SB0 SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M1728 SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Min1 SB1 SubB_0/SR2B_1/Q1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1729 SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Min1 SubB_0/SR2B_1/mux4x1_2/mux2x1_1/Smb SubB_0/SR2B_1/Q1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1730 SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Min1 SubB_0/SR2B_1/mux4x1_2/mux2x1_1/Smb B2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M1731 SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Min1 SB1 B2 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M1732 SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Smb SB0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1733 SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Smb SB0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1734 SubB_0/SR2B_1/mux4x1_2/mux2x1_1/Smb SB1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1735 SubB_0/SR2B_1/mux4x1_2/mux2x1_1/Smb SB1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1736 SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Min2 SB1 SubB_0/SR2B_1/Q1 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M1737 SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Min2 SubB_0/SR2B_1/mux4x1_1/mux2x1_1/Smb SubB_0/SR2B_1/Q1 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M1738 SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Min2 SubB_0/SR2B_1/mux4x1_1/mux2x1_1/Smb SubB_0/SR2B_1/Q2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1739 SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Min2 SB1 SubB_0/SR2B_1/Q2 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1740 SubB_0/SR2B_1/dff3B_1/D SB0 SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M1741 SubB_0/SR2B_1/dff3B_1/D SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Smb SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M1742 SubB_0/SR2B_1/dff3B_1/D SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Smb SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M1743 SubB_0/SR2B_1/dff3B_1/D SB0 SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M1744 SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Min1 SB1 SubB_0/QB0 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1745 SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Min1 SubB_0/SR2B_1/mux4x1_1/mux2x1_1/Smb SubB_0/QB0 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1746 SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Min1 SubB_0/SR2B_1/mux4x1_1/mux2x1_1/Smb B1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M1747 SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Min1 SB1 B1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M1748 SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Smb SB0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1749 SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Smb SB0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1750 SubB_0/SR2B_1/mux4x1_1/mux2x1_1/Smb SB1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1751 SubB_0/SR2B_1/mux4x1_1/mux2x1_1/Smb SB1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1752 SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Min2 SB1 SubB_0/QB0 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M1753 SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Min2 SubB_0/SR2B_1/mux4x1_0/mux2x1_1/Smb SubB_0/QB0 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M1754 SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Min2 SubB_0/SR2B_1/mux4x1_0/mux2x1_1/Smb SubB_0/SR2B_1/Q1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1755 SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Min2 SB1 SubB_0/SR2B_1/Q1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1756 SubB_0/SR2B_1/dff3B_0/D SB0 SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M1757 SubB_0/SR2B_1/dff3B_0/D SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Smb SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M1758 SubB_0/SR2B_1/dff3B_0/D SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Smb SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M1759 SubB_0/SR2B_1/dff3B_0/D SB0 SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M1760 SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Min1 SB1 SR2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M1761 SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Min1 SubB_0/SR2B_1/mux4x1_0/mux2x1_1/Smb SR2 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M1762 SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Min1 SubB_0/SR2B_1/mux4x1_0/mux2x1_1/Smb B0 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M1763 SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Min1 SB1 B0 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M1764 SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Smb SB0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1765 SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Smb SB0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1766 SubB_0/SR2B_1/mux4x1_0/mux2x1_1/Smb SB1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1767 SubB_0/SR2B_1/mux4x1_0/mux2x1_1/Smb SB1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1768 SubB_0/dff3B_0/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1769 SubB_0/dff3B_0/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1770 SubB_0/dff3B_0/gate_0/S SubB_0/dff3B_0/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1771 SubB_0/dff3B_0/gate_0/S SubB_0/dff3B_0/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1772 SubB_0/dff3B_0/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1773 SubB_0/dff3B_0/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1774 nor2_0/in2 SubB_0/dff3B_0/Q Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1775 nor2_0/in2 SubB_0/dff3B_0/Q GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1776 nor2_0/in2 fsm_0/CLK SubB_0/dff3B_0/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1777 nor2_0/in2 SubB_0/dff3B_0/gate_1/S SubB_0/dff3B_0/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1778 SubB_0/dff3B_0/gate_2/Gout SubB_0/dff3B_0/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1779 SubB_0/dff3B_0/gate_2/Gout SubB_0/dff3B_0/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1780 SubB_0/dff3B_0/gate_2/Gout SubB_0/dff3B_0/gate_2/S SubB_0/dff3B_0/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1781 SubB_0/dff3B_0/gate_2/Gout SubB_0/dff3B_0/gate_0/S SubB_0/dff3B_0/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1782 SubB_0/dff3B_0/Qb SubB_0/dff3B_0/Q Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1783 SubB_0/dff3B_0/Qb SubB_0/dff3B_0/Q GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1784 SubB_0/dff3B_0/Q SubB_0/dff3B_0/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1785 SubB_0/dff3B_0/Q SubB_0/dff3B_0/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1786 SubB_0/dff3B_0/gate_3/Gin SubB_0/dff3B_0/gate_1/S SubB_0/dff3B_0/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1787 SubB_0/dff3B_0/gate_3/Gin fsm_0/CLK SubB_0/dff3B_0/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1788 SubB_0/dff3B_0/gate_1/Gin SubB_0/dff3B_0/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1789 SubB_0/dff3B_0/gate_1/Gin SubB_0/dff3B_0/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1790 SubB_0/dff3B_0/gate_2/Gin SubB_0/dff3B_0/gate_0/S SubB_0/dff3B_0/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1791 SubB_0/dff3B_0/gate_2/Gin SubB_0/dff3B_0/gate_2/S SubB_0/dff3B_0/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1792 SubB_0/dff3B_0/gate_0/Gin SubB_0/dff3B_0/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1793 SubB_0/dff3B_0/gate_0/Gin SubB_0/dff3B_0/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1794 SubB_0/dff3B_0/inverter_11/in SubB_0/dff3B_0/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1795 Vdd SubB_0/dff3B_0/D SubB_0/dff3B_0/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1796 SubB_0/dff3B_0/nand2_0/a_n37_n6# SubB_0/dff3B_0/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1797 SubB_0/dff3B_0/inverter_11/in SubB_0/dff3B_0/D SubB_0/dff3B_0/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1798 SubB_0/dff3B_0/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1799 SubB_0/dff3B_0/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1800 Cout SubB_0/xor2_0/nand2_4/nand_in1 Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1801 Vdd SubB_0/xor2_0/nand2_4/nand_in2 Cout Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1802 SubB_0/xor2_0/nand2_4/a_n37_n6# SubB_0/xor2_0/nand2_4/nand_in1 GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1803 Cout SubB_0/xor2_0/nand2_4/nand_in2 SubB_0/xor2_0/nand2_4/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1804 SubB_0/xor2_0/nand2_4/nand_in1 AbS Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1805 Vdd SubB_0/xor2_0/nand2_3/nand_in2 SubB_0/xor2_0/nand2_4/nand_in1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1806 SubB_0/xor2_0/nand2_3/a_n37_n6# AbS GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1807 SubB_0/xor2_0/nand2_4/nand_in1 SubB_0/xor2_0/nand2_3/nand_in2 SubB_0/xor2_0/nand2_3/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1808 SubB_0/xor2_0/nand2_4/nand_in2 SubB_0/xor2_0/nand2_3/nand_in2 Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1809 Vdd SubB_0/dff3B_0/Q SubB_0/xor2_0/nand2_4/nand_in2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1810 SubB_0/xor2_0/nand2_2/a_n37_n6# SubB_0/xor2_0/nand2_3/nand_in2 GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1811 SubB_0/xor2_0/nand2_4/nand_in2 SubB_0/dff3B_0/Q SubB_0/xor2_0/nand2_2/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1812 SubB_0/xor2_0/nand2_3/nand_in2 AbS Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1813 Vdd SubB_0/dff3B_0/Q SubB_0/xor2_0/nand2_3/nand_in2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1814 SubB_0/xor2_0/nand2_1/a_n37_n6# AbS GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1815 SubB_0/xor2_0/nand2_3/nand_in2 SubB_0/dff3B_0/Q SubB_0/xor2_0/nand2_1/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1816 SubB_0/SR2B_0/dff3B_7/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1817 SubB_0/SR2B_0/dff3B_7/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1818 SubB_0/SR2B_0/dff3B_7/gate_0/S SubB_0/SR2B_0/dff3B_7/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1819 SubB_0/SR2B_0/dff3B_7/gate_0/S SubB_0/SR2B_0/dff3B_7/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1820 SubB_0/SR2B_0/dff3B_7/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1821 SubB_0/SR2B_0/dff3B_7/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1822 SubB_0/SR2B_0/dff3B_7/gate_3/Gout SubB_0/SR2B_0/Q7 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1823 SubB_0/SR2B_0/dff3B_7/gate_3/Gout SubB_0/SR2B_0/Q7 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1824 SubB_0/SR2B_0/dff3B_7/gate_3/Gout fsm_0/CLK SubB_0/SR2B_0/dff3B_7/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1825 SubB_0/SR2B_0/dff3B_7/gate_3/Gout SubB_0/SR2B_0/dff3B_7/gate_1/S SubB_0/SR2B_0/dff3B_7/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1826 SubB_0/SR2B_0/dff3B_7/gate_2/Gout SubB_0/SR2B_0/dff3B_7/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1827 SubB_0/SR2B_0/dff3B_7/gate_2/Gout SubB_0/SR2B_0/dff3B_7/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1828 SubB_0/SR2B_0/dff3B_7/gate_2/Gout SubB_0/SR2B_0/dff3B_7/gate_2/S SubB_0/SR2B_0/dff3B_7/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1829 SubB_0/SR2B_0/dff3B_7/gate_2/Gout SubB_0/SR2B_0/dff3B_7/gate_0/S SubB_0/SR2B_0/dff3B_7/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1830 SubB_0/SR2B_0/dff3B_7/Qb SubB_0/SR2B_0/Q7 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1831 SubB_0/SR2B_0/dff3B_7/Qb SubB_0/SR2B_0/Q7 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1832 SubB_0/SR2B_0/Q7 SubB_0/SR2B_0/dff3B_7/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=124p pd=82u as=0p ps=0u 
M1833 SubB_0/SR2B_0/Q7 SubB_0/SR2B_0/dff3B_7/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=75p pd=66u as=0p ps=0u 
M1834 SubB_0/SR2B_0/dff3B_7/gate_3/Gin SubB_0/SR2B_0/dff3B_7/gate_1/S SubB_0/SR2B_0/dff3B_7/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1835 SubB_0/SR2B_0/dff3B_7/gate_3/Gin fsm_0/CLK SubB_0/SR2B_0/dff3B_7/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1836 SubB_0/SR2B_0/dff3B_7/gate_1/Gin SubB_0/SR2B_0/dff3B_7/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1837 SubB_0/SR2B_0/dff3B_7/gate_1/Gin SubB_0/SR2B_0/dff3B_7/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1838 SubB_0/SR2B_0/dff3B_7/gate_2/Gin SubB_0/SR2B_0/dff3B_7/gate_0/S SubB_0/SR2B_0/dff3B_7/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1839 SubB_0/SR2B_0/dff3B_7/gate_2/Gin SubB_0/SR2B_0/dff3B_7/gate_2/S SubB_0/SR2B_0/dff3B_7/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1840 SubB_0/SR2B_0/dff3B_7/gate_0/Gin SubB_0/SR2B_0/dff3B_7/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1841 SubB_0/SR2B_0/dff3B_7/gate_0/Gin SubB_0/SR2B_0/dff3B_7/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1842 SubB_0/SR2B_0/dff3B_7/inverter_11/in SubB_0/SR2B_0/dff3B_7/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1843 Vdd SubB_0/SR2B_0/dff3B_7/D SubB_0/SR2B_0/dff3B_7/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1844 SubB_0/SR2B_0/dff3B_7/nand2_0/a_n37_n6# SubB_0/SR2B_0/dff3B_7/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1845 SubB_0/SR2B_0/dff3B_7/inverter_11/in SubB_0/SR2B_0/dff3B_7/D SubB_0/SR2B_0/dff3B_7/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1846 SubB_0/SR2B_0/dff3B_7/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1847 SubB_0/SR2B_0/dff3B_7/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1848 SubB_0/SR2B_0/dff3B_6/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1849 SubB_0/SR2B_0/dff3B_6/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1850 SubB_0/SR2B_0/dff3B_6/gate_0/S SubB_0/SR2B_0/dff3B_6/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1851 SubB_0/SR2B_0/dff3B_6/gate_0/S SubB_0/SR2B_0/dff3B_6/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1852 SubB_0/SR2B_0/dff3B_6/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1853 SubB_0/SR2B_0/dff3B_6/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1854 SubB_0/SR2B_0/dff3B_6/gate_3/Gout SubB_0/SR2B_0/Q6 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1855 SubB_0/SR2B_0/dff3B_6/gate_3/Gout SubB_0/SR2B_0/Q6 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1856 SubB_0/SR2B_0/dff3B_6/gate_3/Gout fsm_0/CLK SubB_0/SR2B_0/dff3B_6/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1857 SubB_0/SR2B_0/dff3B_6/gate_3/Gout SubB_0/SR2B_0/dff3B_6/gate_1/S SubB_0/SR2B_0/dff3B_6/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1858 SubB_0/SR2B_0/dff3B_6/gate_2/Gout SubB_0/SR2B_0/dff3B_6/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1859 SubB_0/SR2B_0/dff3B_6/gate_2/Gout SubB_0/SR2B_0/dff3B_6/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1860 SubB_0/SR2B_0/dff3B_6/gate_2/Gout SubB_0/SR2B_0/dff3B_6/gate_2/S SubB_0/SR2B_0/dff3B_6/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1861 SubB_0/SR2B_0/dff3B_6/gate_2/Gout SubB_0/SR2B_0/dff3B_6/gate_0/S SubB_0/SR2B_0/dff3B_6/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1862 SubB_0/SR2B_0/dff3B_6/Qb SubB_0/SR2B_0/Q6 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1863 SubB_0/SR2B_0/dff3B_6/Qb SubB_0/SR2B_0/Q6 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1864 SubB_0/SR2B_0/Q6 SubB_0/SR2B_0/dff3B_6/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M1865 SubB_0/SR2B_0/Q6 SubB_0/SR2B_0/dff3B_6/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M1866 SubB_0/SR2B_0/dff3B_6/gate_3/Gin SubB_0/SR2B_0/dff3B_6/gate_1/S SubB_0/SR2B_0/dff3B_6/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1867 SubB_0/SR2B_0/dff3B_6/gate_3/Gin fsm_0/CLK SubB_0/SR2B_0/dff3B_6/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1868 SubB_0/SR2B_0/dff3B_6/gate_1/Gin SubB_0/SR2B_0/dff3B_6/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1869 SubB_0/SR2B_0/dff3B_6/gate_1/Gin SubB_0/SR2B_0/dff3B_6/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1870 SubB_0/SR2B_0/dff3B_6/gate_2/Gin SubB_0/SR2B_0/dff3B_6/gate_0/S SubB_0/SR2B_0/dff3B_6/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1871 SubB_0/SR2B_0/dff3B_6/gate_2/Gin SubB_0/SR2B_0/dff3B_6/gate_2/S SubB_0/SR2B_0/dff3B_6/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1872 SubB_0/SR2B_0/dff3B_6/gate_0/Gin SubB_0/SR2B_0/dff3B_6/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1873 SubB_0/SR2B_0/dff3B_6/gate_0/Gin SubB_0/SR2B_0/dff3B_6/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1874 SubB_0/SR2B_0/dff3B_6/inverter_11/in SubB_0/SR2B_0/dff3B_6/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1875 Vdd SubB_0/SR2B_0/dff3B_6/D SubB_0/SR2B_0/dff3B_6/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1876 SubB_0/SR2B_0/dff3B_6/nand2_0/a_n37_n6# SubB_0/SR2B_0/dff3B_6/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1877 SubB_0/SR2B_0/dff3B_6/inverter_11/in SubB_0/SR2B_0/dff3B_6/D SubB_0/SR2B_0/dff3B_6/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1878 SubB_0/SR2B_0/dff3B_6/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1879 SubB_0/SR2B_0/dff3B_6/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1880 SubB_0/SR2B_0/dff3B_5/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1881 SubB_0/SR2B_0/dff3B_5/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1882 SubB_0/SR2B_0/dff3B_5/gate_0/S SubB_0/SR2B_0/dff3B_5/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1883 SubB_0/SR2B_0/dff3B_5/gate_0/S SubB_0/SR2B_0/dff3B_5/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1884 SubB_0/SR2B_0/dff3B_5/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1885 SubB_0/SR2B_0/dff3B_5/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1886 SubB_0/SR2B_0/dff3B_5/gate_3/Gout SubB_0/SR2B_0/Q5 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1887 SubB_0/SR2B_0/dff3B_5/gate_3/Gout SubB_0/SR2B_0/Q5 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1888 SubB_0/SR2B_0/dff3B_5/gate_3/Gout fsm_0/CLK SubB_0/SR2B_0/dff3B_5/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1889 SubB_0/SR2B_0/dff3B_5/gate_3/Gout SubB_0/SR2B_0/dff3B_5/gate_1/S SubB_0/SR2B_0/dff3B_5/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1890 SubB_0/SR2B_0/dff3B_5/gate_2/Gout SubB_0/SR2B_0/dff3B_5/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1891 SubB_0/SR2B_0/dff3B_5/gate_2/Gout SubB_0/SR2B_0/dff3B_5/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1892 SubB_0/SR2B_0/dff3B_5/gate_2/Gout SubB_0/SR2B_0/dff3B_5/gate_2/S SubB_0/SR2B_0/dff3B_5/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1893 SubB_0/SR2B_0/dff3B_5/gate_2/Gout SubB_0/SR2B_0/dff3B_5/gate_0/S SubB_0/SR2B_0/dff3B_5/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1894 SubB_0/SR2B_0/dff3B_5/Qb SubB_0/SR2B_0/Q5 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1895 SubB_0/SR2B_0/dff3B_5/Qb SubB_0/SR2B_0/Q5 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1896 SubB_0/SR2B_0/Q5 SubB_0/SR2B_0/dff3B_5/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M1897 SubB_0/SR2B_0/Q5 SubB_0/SR2B_0/dff3B_5/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M1898 SubB_0/SR2B_0/dff3B_5/gate_3/Gin SubB_0/SR2B_0/dff3B_5/gate_1/S SubB_0/SR2B_0/dff3B_5/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1899 SubB_0/SR2B_0/dff3B_5/gate_3/Gin fsm_0/CLK SubB_0/SR2B_0/dff3B_5/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1900 SubB_0/SR2B_0/dff3B_5/gate_1/Gin SubB_0/SR2B_0/dff3B_5/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1901 SubB_0/SR2B_0/dff3B_5/gate_1/Gin SubB_0/SR2B_0/dff3B_5/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1902 SubB_0/SR2B_0/dff3B_5/gate_2/Gin SubB_0/SR2B_0/dff3B_5/gate_0/S SubB_0/SR2B_0/dff3B_5/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1903 SubB_0/SR2B_0/dff3B_5/gate_2/Gin SubB_0/SR2B_0/dff3B_5/gate_2/S SubB_0/SR2B_0/dff3B_5/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1904 SubB_0/SR2B_0/dff3B_5/gate_0/Gin SubB_0/SR2B_0/dff3B_5/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1905 SubB_0/SR2B_0/dff3B_5/gate_0/Gin SubB_0/SR2B_0/dff3B_5/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1906 SubB_0/SR2B_0/dff3B_5/inverter_11/in SubB_0/SR2B_0/dff3B_5/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1907 Vdd SubB_0/SR2B_0/dff3B_5/D SubB_0/SR2B_0/dff3B_5/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1908 SubB_0/SR2B_0/dff3B_5/nand2_0/a_n37_n6# SubB_0/SR2B_0/dff3B_5/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1909 SubB_0/SR2B_0/dff3B_5/inverter_11/in SubB_0/SR2B_0/dff3B_5/D SubB_0/SR2B_0/dff3B_5/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1910 SubB_0/SR2B_0/dff3B_5/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1911 SubB_0/SR2B_0/dff3B_5/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1912 SubB_0/SR2B_0/dff3B_4/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1913 SubB_0/SR2B_0/dff3B_4/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1914 SubB_0/SR2B_0/dff3B_4/gate_0/S SubB_0/SR2B_0/dff3B_4/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1915 SubB_0/SR2B_0/dff3B_4/gate_0/S SubB_0/SR2B_0/dff3B_4/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1916 SubB_0/SR2B_0/dff3B_4/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1917 SubB_0/SR2B_0/dff3B_4/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1918 SubB_0/SR2B_0/dff3B_4/gate_3/Gout SubB_0/SR2B_0/Q4 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1919 SubB_0/SR2B_0/dff3B_4/gate_3/Gout SubB_0/SR2B_0/Q4 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1920 SubB_0/SR2B_0/dff3B_4/gate_3/Gout fsm_0/CLK SubB_0/SR2B_0/dff3B_4/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1921 SubB_0/SR2B_0/dff3B_4/gate_3/Gout SubB_0/SR2B_0/dff3B_4/gate_1/S SubB_0/SR2B_0/dff3B_4/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1922 SubB_0/SR2B_0/dff3B_4/gate_2/Gout SubB_0/SR2B_0/dff3B_4/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1923 SubB_0/SR2B_0/dff3B_4/gate_2/Gout SubB_0/SR2B_0/dff3B_4/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1924 SubB_0/SR2B_0/dff3B_4/gate_2/Gout SubB_0/SR2B_0/dff3B_4/gate_2/S SubB_0/SR2B_0/dff3B_4/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1925 SubB_0/SR2B_0/dff3B_4/gate_2/Gout SubB_0/SR2B_0/dff3B_4/gate_0/S SubB_0/SR2B_0/dff3B_4/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1926 SubB_0/SR2B_0/dff3B_4/Qb SubB_0/SR2B_0/Q4 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1927 SubB_0/SR2B_0/dff3B_4/Qb SubB_0/SR2B_0/Q4 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1928 SubB_0/SR2B_0/Q4 SubB_0/SR2B_0/dff3B_4/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M1929 SubB_0/SR2B_0/Q4 SubB_0/SR2B_0/dff3B_4/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M1930 SubB_0/SR2B_0/dff3B_4/gate_3/Gin SubB_0/SR2B_0/dff3B_4/gate_1/S SubB_0/SR2B_0/dff3B_4/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1931 SubB_0/SR2B_0/dff3B_4/gate_3/Gin fsm_0/CLK SubB_0/SR2B_0/dff3B_4/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1932 SubB_0/SR2B_0/dff3B_4/gate_1/Gin SubB_0/SR2B_0/dff3B_4/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1933 SubB_0/SR2B_0/dff3B_4/gate_1/Gin SubB_0/SR2B_0/dff3B_4/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1934 SubB_0/SR2B_0/dff3B_4/gate_2/Gin SubB_0/SR2B_0/dff3B_4/gate_0/S SubB_0/SR2B_0/dff3B_4/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1935 SubB_0/SR2B_0/dff3B_4/gate_2/Gin SubB_0/SR2B_0/dff3B_4/gate_2/S SubB_0/SR2B_0/dff3B_4/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1936 SubB_0/SR2B_0/dff3B_4/gate_0/Gin SubB_0/SR2B_0/dff3B_4/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1937 SubB_0/SR2B_0/dff3B_4/gate_0/Gin SubB_0/SR2B_0/dff3B_4/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1938 SubB_0/SR2B_0/dff3B_4/inverter_11/in SubB_0/SR2B_0/dff3B_4/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1939 Vdd SubB_0/SR2B_0/dff3B_4/D SubB_0/SR2B_0/dff3B_4/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1940 SubB_0/SR2B_0/dff3B_4/nand2_0/a_n37_n6# SubB_0/SR2B_0/dff3B_4/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1941 SubB_0/SR2B_0/dff3B_4/inverter_11/in SubB_0/SR2B_0/dff3B_4/D SubB_0/SR2B_0/dff3B_4/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1942 SubB_0/SR2B_0/dff3B_4/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1943 SubB_0/SR2B_0/dff3B_4/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1944 SubB_0/SR2B_0/dff3B_3/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1945 SubB_0/SR2B_0/dff3B_3/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1946 SubB_0/SR2B_0/dff3B_3/gate_0/S SubB_0/SR2B_0/dff3B_3/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1947 SubB_0/SR2B_0/dff3B_3/gate_0/S SubB_0/SR2B_0/dff3B_3/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1948 SubB_0/SR2B_0/dff3B_3/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1949 SubB_0/SR2B_0/dff3B_3/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1950 SubB_0/SR2B_0/dff3B_3/gate_3/Gout SubB_0/SR2B_0/Q3 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1951 SubB_0/SR2B_0/dff3B_3/gate_3/Gout SubB_0/SR2B_0/Q3 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1952 SubB_0/SR2B_0/dff3B_3/gate_3/Gout fsm_0/CLK SubB_0/SR2B_0/dff3B_3/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1953 SubB_0/SR2B_0/dff3B_3/gate_3/Gout SubB_0/SR2B_0/dff3B_3/gate_1/S SubB_0/SR2B_0/dff3B_3/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1954 SubB_0/SR2B_0/dff3B_3/gate_2/Gout SubB_0/SR2B_0/dff3B_3/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1955 SubB_0/SR2B_0/dff3B_3/gate_2/Gout SubB_0/SR2B_0/dff3B_3/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1956 SubB_0/SR2B_0/dff3B_3/gate_2/Gout SubB_0/SR2B_0/dff3B_3/gate_2/S SubB_0/SR2B_0/dff3B_3/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1957 SubB_0/SR2B_0/dff3B_3/gate_2/Gout SubB_0/SR2B_0/dff3B_3/gate_0/S SubB_0/SR2B_0/dff3B_3/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1958 SubB_0/SR2B_0/dff3B_3/Qb SubB_0/SR2B_0/Q3 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1959 SubB_0/SR2B_0/dff3B_3/Qb SubB_0/SR2B_0/Q3 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1960 SubB_0/SR2B_0/Q3 SubB_0/SR2B_0/dff3B_3/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M1961 SubB_0/SR2B_0/Q3 SubB_0/SR2B_0/dff3B_3/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M1962 SubB_0/SR2B_0/dff3B_3/gate_3/Gin SubB_0/SR2B_0/dff3B_3/gate_1/S SubB_0/SR2B_0/dff3B_3/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1963 SubB_0/SR2B_0/dff3B_3/gate_3/Gin fsm_0/CLK SubB_0/SR2B_0/dff3B_3/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1964 SubB_0/SR2B_0/dff3B_3/gate_1/Gin SubB_0/SR2B_0/dff3B_3/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1965 SubB_0/SR2B_0/dff3B_3/gate_1/Gin SubB_0/SR2B_0/dff3B_3/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1966 SubB_0/SR2B_0/dff3B_3/gate_2/Gin SubB_0/SR2B_0/dff3B_3/gate_0/S SubB_0/SR2B_0/dff3B_3/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1967 SubB_0/SR2B_0/dff3B_3/gate_2/Gin SubB_0/SR2B_0/dff3B_3/gate_2/S SubB_0/SR2B_0/dff3B_3/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1968 SubB_0/SR2B_0/dff3B_3/gate_0/Gin SubB_0/SR2B_0/dff3B_3/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1969 SubB_0/SR2B_0/dff3B_3/gate_0/Gin SubB_0/SR2B_0/dff3B_3/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1970 SubB_0/SR2B_0/dff3B_3/inverter_11/in SubB_0/SR2B_0/dff3B_3/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M1971 Vdd SubB_0/SR2B_0/dff3B_3/D SubB_0/SR2B_0/dff3B_3/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1972 SubB_0/SR2B_0/dff3B_3/nand2_0/a_n37_n6# SubB_0/SR2B_0/dff3B_3/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M1973 SubB_0/SR2B_0/dff3B_3/inverter_11/in SubB_0/SR2B_0/dff3B_3/D SubB_0/SR2B_0/dff3B_3/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1974 SubB_0/SR2B_0/dff3B_3/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1975 SubB_0/SR2B_0/dff3B_3/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1976 SubB_0/SR2B_0/dff3B_2/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1977 SubB_0/SR2B_0/dff3B_2/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1978 SubB_0/SR2B_0/dff3B_2/gate_0/S SubB_0/SR2B_0/dff3B_2/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1979 SubB_0/SR2B_0/dff3B_2/gate_0/S SubB_0/SR2B_0/dff3B_2/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1980 SubB_0/SR2B_0/dff3B_2/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1981 SubB_0/SR2B_0/dff3B_2/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1982 SubB_0/SR2B_0/dff3B_2/gate_3/Gout SubB_0/SR2B_0/Q2 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1983 SubB_0/SR2B_0/dff3B_2/gate_3/Gout SubB_0/SR2B_0/Q2 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1984 SubB_0/SR2B_0/dff3B_2/gate_3/Gout fsm_0/CLK SubB_0/SR2B_0/dff3B_2/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1985 SubB_0/SR2B_0/dff3B_2/gate_3/Gout SubB_0/SR2B_0/dff3B_2/gate_1/S SubB_0/SR2B_0/dff3B_2/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1986 SubB_0/SR2B_0/dff3B_2/gate_2/Gout SubB_0/SR2B_0/dff3B_2/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M1987 SubB_0/SR2B_0/dff3B_2/gate_2/Gout SubB_0/SR2B_0/dff3B_2/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M1988 SubB_0/SR2B_0/dff3B_2/gate_2/Gout SubB_0/SR2B_0/dff3B_2/gate_2/S SubB_0/SR2B_0/dff3B_2/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M1989 SubB_0/SR2B_0/dff3B_2/gate_2/Gout SubB_0/SR2B_0/dff3B_2/gate_0/S SubB_0/SR2B_0/dff3B_2/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M1990 SubB_0/SR2B_0/dff3B_2/Qb SubB_0/SR2B_0/Q2 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M1991 SubB_0/SR2B_0/dff3B_2/Qb SubB_0/SR2B_0/Q2 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M1992 SubB_0/SR2B_0/Q2 SubB_0/SR2B_0/dff3B_2/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M1993 SubB_0/SR2B_0/Q2 SubB_0/SR2B_0/dff3B_2/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M1994 SubB_0/SR2B_0/dff3B_2/gate_3/Gin SubB_0/SR2B_0/dff3B_2/gate_1/S SubB_0/SR2B_0/dff3B_2/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1995 SubB_0/SR2B_0/dff3B_2/gate_3/Gin fsm_0/CLK SubB_0/SR2B_0/dff3B_2/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M1996 SubB_0/SR2B_0/dff3B_2/gate_1/Gin SubB_0/SR2B_0/dff3B_2/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1997 SubB_0/SR2B_0/dff3B_2/gate_1/Gin SubB_0/SR2B_0/dff3B_2/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1998 SubB_0/SR2B_0/dff3B_2/gate_2/Gin SubB_0/SR2B_0/dff3B_2/gate_0/S SubB_0/SR2B_0/dff3B_2/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M1999 SubB_0/SR2B_0/dff3B_2/gate_2/Gin SubB_0/SR2B_0/dff3B_2/gate_2/S SubB_0/SR2B_0/dff3B_2/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2000 SubB_0/SR2B_0/dff3B_2/gate_0/Gin SubB_0/SR2B_0/dff3B_2/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2001 SubB_0/SR2B_0/dff3B_2/gate_0/Gin SubB_0/SR2B_0/dff3B_2/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2002 SubB_0/SR2B_0/dff3B_2/inverter_11/in SubB_0/SR2B_0/dff3B_2/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2003 Vdd SubB_0/SR2B_0/dff3B_2/D SubB_0/SR2B_0/dff3B_2/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2004 SubB_0/SR2B_0/dff3B_2/nand2_0/a_n37_n6# SubB_0/SR2B_0/dff3B_2/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2005 SubB_0/SR2B_0/dff3B_2/inverter_11/in SubB_0/SR2B_0/dff3B_2/D SubB_0/SR2B_0/dff3B_2/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2006 SubB_0/SR2B_0/dff3B_2/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2007 SubB_0/SR2B_0/dff3B_2/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2008 SubB_0/SR2B_0/dff3B_1/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2009 SubB_0/SR2B_0/dff3B_1/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2010 SubB_0/SR2B_0/dff3B_1/gate_0/S SubB_0/SR2B_0/dff3B_1/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2011 SubB_0/SR2B_0/dff3B_1/gate_0/S SubB_0/SR2B_0/dff3B_1/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2012 SubB_0/SR2B_0/dff3B_1/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2013 SubB_0/SR2B_0/dff3B_1/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2014 SubB_0/SR2B_0/dff3B_1/gate_3/Gout SubB_0/SR2B_0/Q1 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2015 SubB_0/SR2B_0/dff3B_1/gate_3/Gout SubB_0/SR2B_0/Q1 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2016 SubB_0/SR2B_0/dff3B_1/gate_3/Gout fsm_0/CLK SubB_0/SR2B_0/dff3B_1/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2017 SubB_0/SR2B_0/dff3B_1/gate_3/Gout SubB_0/SR2B_0/dff3B_1/gate_1/S SubB_0/SR2B_0/dff3B_1/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2018 SubB_0/SR2B_0/dff3B_1/gate_2/Gout SubB_0/SR2B_0/dff3B_1/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2019 SubB_0/SR2B_0/dff3B_1/gate_2/Gout SubB_0/SR2B_0/dff3B_1/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2020 SubB_0/SR2B_0/dff3B_1/gate_2/Gout SubB_0/SR2B_0/dff3B_1/gate_2/S SubB_0/SR2B_0/dff3B_1/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2021 SubB_0/SR2B_0/dff3B_1/gate_2/Gout SubB_0/SR2B_0/dff3B_1/gate_0/S SubB_0/SR2B_0/dff3B_1/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2022 SubB_0/SR2B_0/dff3B_1/Qb SubB_0/SR2B_0/Q1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2023 SubB_0/SR2B_0/dff3B_1/Qb SubB_0/SR2B_0/Q1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2024 SubB_0/SR2B_0/Q1 SubB_0/SR2B_0/dff3B_1/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M2025 SubB_0/SR2B_0/Q1 SubB_0/SR2B_0/dff3B_1/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M2026 SubB_0/SR2B_0/dff3B_1/gate_3/Gin SubB_0/SR2B_0/dff3B_1/gate_1/S SubB_0/SR2B_0/dff3B_1/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2027 SubB_0/SR2B_0/dff3B_1/gate_3/Gin fsm_0/CLK SubB_0/SR2B_0/dff3B_1/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2028 SubB_0/SR2B_0/dff3B_1/gate_1/Gin SubB_0/SR2B_0/dff3B_1/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2029 SubB_0/SR2B_0/dff3B_1/gate_1/Gin SubB_0/SR2B_0/dff3B_1/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2030 SubB_0/SR2B_0/dff3B_1/gate_2/Gin SubB_0/SR2B_0/dff3B_1/gate_0/S SubB_0/SR2B_0/dff3B_1/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2031 SubB_0/SR2B_0/dff3B_1/gate_2/Gin SubB_0/SR2B_0/dff3B_1/gate_2/S SubB_0/SR2B_0/dff3B_1/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2032 SubB_0/SR2B_0/dff3B_1/gate_0/Gin SubB_0/SR2B_0/dff3B_1/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2033 SubB_0/SR2B_0/dff3B_1/gate_0/Gin SubB_0/SR2B_0/dff3B_1/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2034 SubB_0/SR2B_0/dff3B_1/inverter_11/in SubB_0/SR2B_0/dff3B_1/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2035 Vdd SubB_0/SR2B_0/dff3B_1/D SubB_0/SR2B_0/dff3B_1/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2036 SubB_0/SR2B_0/dff3B_1/nand2_0/a_n37_n6# SubB_0/SR2B_0/dff3B_1/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2037 SubB_0/SR2B_0/dff3B_1/inverter_11/in SubB_0/SR2B_0/dff3B_1/D SubB_0/SR2B_0/dff3B_1/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2038 SubB_0/SR2B_0/dff3B_1/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2039 SubB_0/SR2B_0/dff3B_1/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2040 SubB_0/SR2B_0/dff3B_0/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2041 SubB_0/SR2B_0/dff3B_0/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2042 SubB_0/SR2B_0/dff3B_0/gate_0/S SubB_0/SR2B_0/dff3B_0/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2043 SubB_0/SR2B_0/dff3B_0/gate_0/S SubB_0/SR2B_0/dff3B_0/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2044 SubB_0/SR2B_0/dff3B_0/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2045 SubB_0/SR2B_0/dff3B_0/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2046 SubB_0/SR2B_0/dff3B_0/gate_3/Gout SubB_0/QA0 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2047 SubB_0/SR2B_0/dff3B_0/gate_3/Gout SubB_0/QA0 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2048 SubB_0/SR2B_0/dff3B_0/gate_3/Gout fsm_0/CLK SubB_0/SR2B_0/dff3B_0/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2049 SubB_0/SR2B_0/dff3B_0/gate_3/Gout SubB_0/SR2B_0/dff3B_0/gate_1/S SubB_0/SR2B_0/dff3B_0/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2050 SubB_0/SR2B_0/dff3B_0/gate_2/Gout SubB_0/SR2B_0/dff3B_0/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2051 SubB_0/SR2B_0/dff3B_0/gate_2/Gout SubB_0/SR2B_0/dff3B_0/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2052 SubB_0/SR2B_0/dff3B_0/gate_2/Gout SubB_0/SR2B_0/dff3B_0/gate_2/S SubB_0/SR2B_0/dff3B_0/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2053 SubB_0/SR2B_0/dff3B_0/gate_2/Gout SubB_0/SR2B_0/dff3B_0/gate_0/S SubB_0/SR2B_0/dff3B_0/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2054 SubB_0/SR2B_0/dff3B_0/Qb SubB_0/QA0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2055 SubB_0/SR2B_0/dff3B_0/Qb SubB_0/QA0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2056 SubB_0/QA0 SubB_0/SR2B_0/dff3B_0/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=173p pd=112u as=0p ps=0u 
M2057 SubB_0/QA0 SubB_0/SR2B_0/dff3B_0/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=103p pd=90u as=0p ps=0u 
M2058 SubB_0/SR2B_0/dff3B_0/gate_3/Gin SubB_0/SR2B_0/dff3B_0/gate_1/S SubB_0/SR2B_0/dff3B_0/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2059 SubB_0/SR2B_0/dff3B_0/gate_3/Gin fsm_0/CLK SubB_0/SR2B_0/dff3B_0/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2060 SubB_0/SR2B_0/dff3B_0/gate_1/Gin SubB_0/SR2B_0/dff3B_0/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2061 SubB_0/SR2B_0/dff3B_0/gate_1/Gin SubB_0/SR2B_0/dff3B_0/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2062 SubB_0/SR2B_0/dff3B_0/gate_2/Gin SubB_0/SR2B_0/dff3B_0/gate_0/S SubB_0/SR2B_0/dff3B_0/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2063 SubB_0/SR2B_0/dff3B_0/gate_2/Gin SubB_0/SR2B_0/dff3B_0/gate_2/S SubB_0/SR2B_0/dff3B_0/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2064 SubB_0/SR2B_0/dff3B_0/gate_0/Gin SubB_0/SR2B_0/dff3B_0/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2065 SubB_0/SR2B_0/dff3B_0/gate_0/Gin SubB_0/SR2B_0/dff3B_0/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2066 SubB_0/SR2B_0/dff3B_0/inverter_11/in SubB_0/SR2B_0/dff3B_0/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2067 Vdd SubB_0/SR2B_0/dff3B_0/D SubB_0/SR2B_0/dff3B_0/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2068 SubB_0/SR2B_0/dff3B_0/nand2_0/a_n37_n6# SubB_0/SR2B_0/dff3B_0/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2069 SubB_0/SR2B_0/dff3B_0/inverter_11/in SubB_0/SR2B_0/dff3B_0/D SubB_0/SR2B_0/dff3B_0/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2070 SubB_0/SR2B_0/dff3B_0/inverter_7/out fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2071 SubB_0/SR2B_0/dff3B_0/inverter_7/out fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2072 SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Min2 SA1 SubB_0/SR2B_0/Q7 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M2073 SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Min2 SubB_0/SR2B_0/mux4x1_7/mux2x1_1/Smb SubB_0/SR2B_0/Q7 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M2074 SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Min2 SubB_0/SR2B_0/mux4x1_7/mux2x1_1/Smb SubB_0/QA0 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2075 SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Min2 SA1 SubB_0/QA0 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2076 SubB_0/SR2B_0/dff3B_7/D SA0 SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M2077 SubB_0/SR2B_0/dff3B_7/D SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Smb SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M2078 SubB_0/SR2B_0/dff3B_7/D SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Smb SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M2079 SubB_0/SR2B_0/dff3B_7/D SA0 SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M2080 SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Min1 SA1 SubB_0/SR2B_0/Q6 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2081 SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Min1 SubB_0/SR2B_0/mux4x1_7/mux2x1_1/Smb SubB_0/SR2B_0/Q6 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2082 SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Min1 SubB_0/SR2B_0/mux4x1_7/mux2x1_1/Smb A7 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M2083 SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Min1 SA1 A7 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M2084 SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Smb SA0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2085 SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Smb SA0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2086 SubB_0/SR2B_0/mux4x1_7/mux2x1_1/Smb SA1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2087 SubB_0/SR2B_0/mux4x1_7/mux2x1_1/Smb SA1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2088 SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Min2 SA1 SubB_0/SR2B_0/Q6 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M2089 SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Min2 SubB_0/SR2B_0/mux4x1_6/mux2x1_1/Smb SubB_0/SR2B_0/Q6 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M2090 SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Min2 SubB_0/SR2B_0/mux4x1_6/mux2x1_1/Smb SubB_0/SR2B_0/Q7 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2091 SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Min2 SA1 SubB_0/SR2B_0/Q7 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2092 SubB_0/SR2B_0/dff3B_6/D SA0 SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M2093 SubB_0/SR2B_0/dff3B_6/D SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Smb SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M2094 SubB_0/SR2B_0/dff3B_6/D SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Smb SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M2095 SubB_0/SR2B_0/dff3B_6/D SA0 SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M2096 SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Min1 SA1 SubB_0/SR2B_0/Q5 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2097 SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Min1 SubB_0/SR2B_0/mux4x1_6/mux2x1_1/Smb SubB_0/SR2B_0/Q5 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2098 SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Min1 SubB_0/SR2B_0/mux4x1_6/mux2x1_1/Smb A6 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M2099 SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Min1 SA1 A6 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M2100 SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Smb SA0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2101 SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Smb SA0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2102 SubB_0/SR2B_0/mux4x1_6/mux2x1_1/Smb SA1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2103 SubB_0/SR2B_0/mux4x1_6/mux2x1_1/Smb SA1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2104 SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Min2 SA1 SubB_0/SR2B_0/Q5 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M2105 SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Min2 SubB_0/SR2B_0/mux4x1_5/mux2x1_1/Smb SubB_0/SR2B_0/Q5 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M2106 SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Min2 SubB_0/SR2B_0/mux4x1_5/mux2x1_1/Smb SubB_0/SR2B_0/Q6 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2107 SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Min2 SA1 SubB_0/SR2B_0/Q6 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2108 SubB_0/SR2B_0/dff3B_5/D SA0 SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M2109 SubB_0/SR2B_0/dff3B_5/D SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Smb SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M2110 SubB_0/SR2B_0/dff3B_5/D SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Smb SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M2111 SubB_0/SR2B_0/dff3B_5/D SA0 SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M2112 SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Min1 SA1 SubB_0/SR2B_0/Q4 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2113 SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Min1 SubB_0/SR2B_0/mux4x1_5/mux2x1_1/Smb SubB_0/SR2B_0/Q4 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2114 SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Min1 SubB_0/SR2B_0/mux4x1_5/mux2x1_1/Smb A5 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M2115 SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Min1 SA1 A5 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M2116 SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Smb SA0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2117 SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Smb SA0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2118 SubB_0/SR2B_0/mux4x1_5/mux2x1_1/Smb SA1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2119 SubB_0/SR2B_0/mux4x1_5/mux2x1_1/Smb SA1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2120 SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Min2 SA1 SubB_0/SR2B_0/Q4 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M2121 SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Min2 SubB_0/SR2B_0/mux4x1_4/mux2x1_1/Smb SubB_0/SR2B_0/Q4 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M2122 SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Min2 SubB_0/SR2B_0/mux4x1_4/mux2x1_1/Smb SubB_0/SR2B_0/Q5 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2123 SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Min2 SA1 SubB_0/SR2B_0/Q5 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2124 SubB_0/SR2B_0/dff3B_4/D SA0 SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M2125 SubB_0/SR2B_0/dff3B_4/D SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Smb SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M2126 SubB_0/SR2B_0/dff3B_4/D SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Smb SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M2127 SubB_0/SR2B_0/dff3B_4/D SA0 SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M2128 SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Min1 SA1 SubB_0/SR2B_0/Q3 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2129 SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Min1 SubB_0/SR2B_0/mux4x1_4/mux2x1_1/Smb SubB_0/SR2B_0/Q3 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2130 SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Min1 SubB_0/SR2B_0/mux4x1_4/mux2x1_1/Smb A4 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M2131 SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Min1 SA1 A4 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M2132 SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Smb SA0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2133 SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Smb SA0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2134 SubB_0/SR2B_0/mux4x1_4/mux2x1_1/Smb SA1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2135 SubB_0/SR2B_0/mux4x1_4/mux2x1_1/Smb SA1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2136 SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Min2 SA1 SubB_0/SR2B_0/Q3 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M2137 SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Min2 SubB_0/SR2B_0/mux4x1_3/mux2x1_1/Smb SubB_0/SR2B_0/Q3 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M2138 SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Min2 SubB_0/SR2B_0/mux4x1_3/mux2x1_1/Smb SubB_0/SR2B_0/Q4 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2139 SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Min2 SA1 SubB_0/SR2B_0/Q4 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2140 SubB_0/SR2B_0/dff3B_3/D SA0 SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M2141 SubB_0/SR2B_0/dff3B_3/D SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Smb SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M2142 SubB_0/SR2B_0/dff3B_3/D SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Smb SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M2143 SubB_0/SR2B_0/dff3B_3/D SA0 SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M2144 SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Min1 SA1 SubB_0/SR2B_0/Q2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2145 SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Min1 SubB_0/SR2B_0/mux4x1_3/mux2x1_1/Smb SubB_0/SR2B_0/Q2 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2146 SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Min1 SubB_0/SR2B_0/mux4x1_3/mux2x1_1/Smb A3 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M2147 SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Min1 SA1 A3 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M2148 SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Smb SA0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2149 SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Smb SA0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2150 SubB_0/SR2B_0/mux4x1_3/mux2x1_1/Smb SA1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2151 SubB_0/SR2B_0/mux4x1_3/mux2x1_1/Smb SA1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2152 SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Min2 SA1 SubB_0/SR2B_0/Q2 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M2153 SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Min2 SubB_0/SR2B_0/mux4x1_2/mux2x1_1/Smb SubB_0/SR2B_0/Q2 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M2154 SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Min2 SubB_0/SR2B_0/mux4x1_2/mux2x1_1/Smb SubB_0/SR2B_0/Q3 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2155 SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Min2 SA1 SubB_0/SR2B_0/Q3 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2156 SubB_0/SR2B_0/dff3B_2/D SA0 SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M2157 SubB_0/SR2B_0/dff3B_2/D SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Smb SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M2158 SubB_0/SR2B_0/dff3B_2/D SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Smb SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M2159 SubB_0/SR2B_0/dff3B_2/D SA0 SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M2160 SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Min1 SA1 SubB_0/SR2B_0/Q1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2161 SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Min1 SubB_0/SR2B_0/mux4x1_2/mux2x1_1/Smb SubB_0/SR2B_0/Q1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2162 SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Min1 SubB_0/SR2B_0/mux4x1_2/mux2x1_1/Smb A2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M2163 SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Min1 SA1 A2 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M2164 SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Smb SA0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2165 SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Smb SA0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2166 SubB_0/SR2B_0/mux4x1_2/mux2x1_1/Smb SA1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2167 SubB_0/SR2B_0/mux4x1_2/mux2x1_1/Smb SA1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2168 SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Min2 SA1 SubB_0/SR2B_0/Q1 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M2169 SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Min2 SubB_0/SR2B_0/mux4x1_1/mux2x1_1/Smb SubB_0/SR2B_0/Q1 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M2170 SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Min2 SubB_0/SR2B_0/mux4x1_1/mux2x1_1/Smb SubB_0/SR2B_0/Q2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2171 SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Min2 SA1 SubB_0/SR2B_0/Q2 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2172 SubB_0/SR2B_0/dff3B_1/D SA0 SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M2173 SubB_0/SR2B_0/dff3B_1/D SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Smb SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M2174 SubB_0/SR2B_0/dff3B_1/D SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Smb SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M2175 SubB_0/SR2B_0/dff3B_1/D SA0 SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M2176 SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Min1 SA1 SubB_0/QA0 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2177 SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Min1 SubB_0/SR2B_0/mux4x1_1/mux2x1_1/Smb SubB_0/QA0 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2178 SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Min1 SubB_0/SR2B_0/mux4x1_1/mux2x1_1/Smb A1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M2179 SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Min1 SA1 A1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M2180 SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Smb SA0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2181 SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Smb SA0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2182 SubB_0/SR2B_0/mux4x1_1/mux2x1_1/Smb SA1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2183 SubB_0/SR2B_0/mux4x1_1/mux2x1_1/Smb SA1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2184 SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Min2 SA1 SubB_0/QA0 Vdd pfet w=6u l=2u
+ ad=147p pd=90u as=0p ps=0u 
M2185 SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Min2 SubB_0/SR2B_0/mux4x1_0/mux2x1_1/Smb SubB_0/QA0 Gnd nfet w=3u l=2u
+ ad=84p pd=72u as=0p ps=0u 
M2186 SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Min2 SubB_0/SR2B_0/mux4x1_0/mux2x1_1/Smb SubB_0/SR2B_0/Q1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2187 SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Min2 SA1 SubB_0/SR2B_0/Q1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2188 SubB_0/SR2B_0/dff3B_0/D SA0 SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Min2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M2189 SubB_0/SR2B_0/dff3B_0/D SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Smb SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Min2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M2190 SubB_0/SR2B_0/dff3B_0/D SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Smb SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Min1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=147p ps=90u 
M2191 SubB_0/SR2B_0/dff3B_0/D SA0 SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Min1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=84p ps=72u 
M2192 SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Min1 SA1 SR Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M2193 SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Min1 SubB_0/SR2B_0/mux4x1_0/mux2x1_1/Smb SR Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M2194 SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Min1 SubB_0/SR2B_0/mux4x1_0/mux2x1_1/Smb A0 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=49p ps=30u 
M2195 SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Min1 SA1 A0 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=28p ps=24u 
M2196 SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Smb SA0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2197 SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Smb SA0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2198 SubB_0/SR2B_0/mux4x1_0/mux2x1_1/Smb SA1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2199 SubB_0/SR2B_0/mux4x1_0/mux2x1_1/Smb SA1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2200 SubB_0/dff3B_0/D SubB_0/abs_0/nor2_0/out Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2201 SubB_0/dff3B_0/D SubB_0/abs_0/nor2_0/out GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2202 SubB_0/abs_0/nor2_0/a_n37_6# SubB_0/abs_0/nor2_0/in1 Vdd Vdd pfet w=6u l=2u
+ ad=12p pd=16u as=0p ps=0u 
M2203 SubB_0/abs_0/nor2_0/out SubB_0/abs_0/nor2_0/in2 SubB_0/abs_0/nor2_0/a_n37_6# Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2204 SubB_0/abs_0/nor2_0/out SubB_0/abs_0/nor2_0/in1 GND Gnd nfet w=3u l=2u
+ ad=22p pd=20u as=0p ps=0u 
M2205 GND SubB_0/abs_0/nor2_0/in2 SubB_0/abs_0/nor2_0/out Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2206 SubB_0/abs_0/sum SubB_0/abs_0/ha_1/xor2_0/nand2_4/nand_in1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2207 Vdd SubB_0/abs_0/ha_1/xor2_0/nand2_4/nand_in2 SubB_0/abs_0/sum Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2208 SubB_0/abs_0/ha_1/xor2_0/nand2_4/a_n37_n6# SubB_0/abs_0/ha_1/xor2_0/nand2_4/nand_in1 GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2209 SubB_0/abs_0/sum SubB_0/abs_0/ha_1/xor2_0/nand2_4/nand_in2 SubB_0/abs_0/ha_1/xor2_0/nand2_4/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2210 SubB_0/abs_0/ha_1/xor2_0/nand2_4/nand_in1 SubB_0/abs_0/ha_1/ha_in1 Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2211 Vdd SubB_0/abs_0/ha_1/xor2_0/nand2_3/nand_in2 SubB_0/abs_0/ha_1/xor2_0/nand2_4/nand_in1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2212 SubB_0/abs_0/ha_1/xor2_0/nand2_3/a_n37_n6# SubB_0/abs_0/ha_1/ha_in1 GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2213 SubB_0/abs_0/ha_1/xor2_0/nand2_4/nand_in1 SubB_0/abs_0/ha_1/xor2_0/nand2_3/nand_in2 SubB_0/abs_0/ha_1/xor2_0/nand2_3/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2214 SubB_0/abs_0/ha_1/xor2_0/nand2_4/nand_in2 SubB_0/abs_0/ha_1/xor2_0/nand2_3/nand_in2 Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2215 Vdd SubB_0/abs_0/cin SubB_0/abs_0/ha_1/xor2_0/nand2_4/nand_in2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2216 SubB_0/abs_0/ha_1/xor2_0/nand2_2/a_n37_n6# SubB_0/abs_0/ha_1/xor2_0/nand2_3/nand_in2 GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2217 SubB_0/abs_0/ha_1/xor2_0/nand2_4/nand_in2 SubB_0/abs_0/cin SubB_0/abs_0/ha_1/xor2_0/nand2_2/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2218 SubB_0/abs_0/ha_1/xor2_0/nand2_3/nand_in2 SubB_0/abs_0/ha_1/ha_in1 Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2219 Vdd SubB_0/abs_0/cin SubB_0/abs_0/ha_1/xor2_0/nand2_3/nand_in2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2220 SubB_0/abs_0/ha_1/xor2_0/nand2_1/a_n37_n6# SubB_0/abs_0/ha_1/ha_in1 GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2221 SubB_0/abs_0/ha_1/xor2_0/nand2_3/nand_in2 SubB_0/abs_0/cin SubB_0/abs_0/ha_1/xor2_0/nand2_1/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2222 SubB_0/abs_0/nor2_0/in2 SubB_0/abs_0/ha_1/not1_0/not_in Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2223 SubB_0/abs_0/nor2_0/in2 SubB_0/abs_0/ha_1/not1_0/not_in GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2224 SubB_0/abs_0/ha_1/not1_0/not_in SubB_0/abs_0/ha_1/ha_in1 Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2225 Vdd SubB_0/abs_0/cin SubB_0/abs_0/ha_1/not1_0/not_in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2226 SubB_0/abs_0/ha_1/nand2_0/a_n37_n6# SubB_0/abs_0/ha_1/ha_in1 GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2227 SubB_0/abs_0/ha_1/not1_0/not_in SubB_0/abs_0/cin SubB_0/abs_0/ha_1/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2228 SubB_0/abs_0/ha_1/ha_in1 SubB_0/abs_0/ha_0/xor2_0/nand2_4/nand_in1 Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2229 Vdd SubB_0/abs_0/ha_0/xor2_0/nand2_4/nand_in2 SubB_0/abs_0/ha_1/ha_in1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2230 SubB_0/abs_0/ha_0/xor2_0/nand2_4/a_n37_n6# SubB_0/abs_0/ha_0/xor2_0/nand2_4/nand_in1 GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2231 SubB_0/abs_0/ha_1/ha_in1 SubB_0/abs_0/ha_0/xor2_0/nand2_4/nand_in2 SubB_0/abs_0/ha_0/xor2_0/nand2_4/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2232 SubB_0/abs_0/ha_0/xor2_0/nand2_4/nand_in1 SubB_0/QA0 Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2233 Vdd SubB_0/abs_0/ha_0/xor2_0/nand2_3/nand_in2 SubB_0/abs_0/ha_0/xor2_0/nand2_4/nand_in1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2234 SubB_0/abs_0/ha_0/xor2_0/nand2_3/a_n37_n6# SubB_0/QA0 GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2235 SubB_0/abs_0/ha_0/xor2_0/nand2_4/nand_in1 SubB_0/abs_0/ha_0/xor2_0/nand2_3/nand_in2 SubB_0/abs_0/ha_0/xor2_0/nand2_3/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2236 SubB_0/abs_0/ha_0/xor2_0/nand2_4/nand_in2 SubB_0/abs_0/ha_0/xor2_0/nand2_3/nand_in2 Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2237 Vdd SubB_0/abs_0/ha_0/ha_in2 SubB_0/abs_0/ha_0/xor2_0/nand2_4/nand_in2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2238 SubB_0/abs_0/ha_0/xor2_0/nand2_2/a_n37_n6# SubB_0/abs_0/ha_0/xor2_0/nand2_3/nand_in2 GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2239 SubB_0/abs_0/ha_0/xor2_0/nand2_4/nand_in2 SubB_0/abs_0/ha_0/ha_in2 SubB_0/abs_0/ha_0/xor2_0/nand2_2/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2240 SubB_0/abs_0/ha_0/xor2_0/nand2_3/nand_in2 SubB_0/QA0 Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2241 Vdd SubB_0/abs_0/ha_0/ha_in2 SubB_0/abs_0/ha_0/xor2_0/nand2_3/nand_in2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2242 SubB_0/abs_0/ha_0/xor2_0/nand2_1/a_n37_n6# SubB_0/QA0 GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2243 SubB_0/abs_0/ha_0/xor2_0/nand2_3/nand_in2 SubB_0/abs_0/ha_0/ha_in2 SubB_0/abs_0/ha_0/xor2_0/nand2_1/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2244 SubB_0/abs_0/nor2_0/in1 SubB_0/abs_0/ha_0/not1_0/not_in Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2245 SubB_0/abs_0/nor2_0/in1 SubB_0/abs_0/ha_0/not1_0/not_in GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2246 SubB_0/abs_0/ha_0/not1_0/not_in SubB_0/QA0 Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2247 Vdd SubB_0/abs_0/ha_0/ha_in2 SubB_0/abs_0/ha_0/not1_0/not_in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2248 SubB_0/abs_0/ha_0/nand2_0/a_n37_n6# SubB_0/QA0 GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2249 SubB_0/abs_0/ha_0/not1_0/not_in SubB_0/abs_0/ha_0/ha_in2 SubB_0/abs_0/ha_0/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2250 SubB_0/abs_0/ha_0/ha_in2 SubB_0/abs_0/xor2_0/nand2_4/nand_in1 Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2251 Vdd SubB_0/abs_0/xor2_0/nand2_4/nand_in2 SubB_0/abs_0/ha_0/ha_in2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2252 SubB_0/abs_0/xor2_0/nand2_4/a_n37_n6# SubB_0/abs_0/xor2_0/nand2_4/nand_in1 GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2253 SubB_0/abs_0/ha_0/ha_in2 SubB_0/abs_0/xor2_0/nand2_4/nand_in2 SubB_0/abs_0/xor2_0/nand2_4/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2254 SubB_0/abs_0/xor2_0/nand2_4/nand_in1 AbS Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2255 Vdd SubB_0/abs_0/xor2_0/nand2_3/nand_in2 SubB_0/abs_0/xor2_0/nand2_4/nand_in1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2256 SubB_0/abs_0/xor2_0/nand2_3/a_n37_n6# AbS GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2257 SubB_0/abs_0/xor2_0/nand2_4/nand_in1 SubB_0/abs_0/xor2_0/nand2_3/nand_in2 SubB_0/abs_0/xor2_0/nand2_3/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2258 SubB_0/abs_0/xor2_0/nand2_4/nand_in2 SubB_0/abs_0/xor2_0/nand2_3/nand_in2 Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2259 Vdd SubB_0/QB0 SubB_0/abs_0/xor2_0/nand2_4/nand_in2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2260 SubB_0/abs_0/xor2_0/nand2_2/a_n37_n6# SubB_0/abs_0/xor2_0/nand2_3/nand_in2 GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2261 SubB_0/abs_0/xor2_0/nand2_4/nand_in2 SubB_0/QB0 SubB_0/abs_0/xor2_0/nand2_2/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2262 SubB_0/abs_0/xor2_0/nand2_3/nand_in2 AbS Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2263 Vdd SubB_0/QB0 SubB_0/abs_0/xor2_0/nand2_3/nand_in2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2264 SubB_0/abs_0/xor2_0/nand2_1/a_n37_n6# AbS GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2265 SubB_0/abs_0/xor2_0/nand2_3/nand_in2 SubB_0/QB0 SubB_0/abs_0/xor2_0/nand2_1/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2266 SubB_0/abs_0/cin SubB_0/mux2x1_0/Sm AbS Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=49p ps=30u 
M2267 SubB_0/abs_0/cin fsm_0/A3 AbS Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=28p ps=24u 
M2268 SubB_0/abs_0/cin fsm_0/A3 SubB_0/dff3B_0/Q Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2269 SubB_0/abs_0/cin SubB_0/mux2x1_0/Sm SubB_0/dff3B_0/Q Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2270 SubB_0/mux2x1_0/Sm fsm_0/A3 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2271 SubB_0/mux2x1_0/Sm fsm_0/A3 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2272 nor2_0/a_n37_6# nor2_0/in1 Vdd Vdd pfet w=6u l=2u
+ ad=12p pd=16u as=0p ps=0u 
M2273 nor2_0/out nor2_0/in2 nor2_0/a_n37_6# Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2274 nor2_0/out nor2_0/in1 GND Gnd nfet w=3u l=2u
+ ad=22p pd=20u as=0p ps=0u 
M2275 GND nor2_0/in2 nor2_0/out Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2276 nor2_0/in1 nor2_0/in2 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2277 nor2_0/in1 nor2_0/in2 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2278 SB1 fsm_0/nor2_3/out Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2279 SB1 fsm_0/nor2_3/out GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2280 SA1 fsm_0/nor2_4/out Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2281 SA1 fsm_0/nor2_4/out GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2282 SS0 fsm_0/inverter_9/in Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2283 SS0 fsm_0/inverter_9/in GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2284 fsm_0/nor2_3/a_n37_6# SS0 Vdd Vdd pfet w=6u l=2u
+ ad=12p pd=16u as=0p ps=0u 
M2285 fsm_0/nor2_3/out SB0 fsm_0/nor2_3/a_n37_6# Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2286 fsm_0/nor2_3/out SS0 GND Gnd nfet w=3u l=2u
+ ad=22p pd=20u as=0p ps=0u 
M2287 GND SB0 fsm_0/nor2_3/out Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2288 SB0 fsm_0/inverter_8/in Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2289 SB0 fsm_0/inverter_8/in GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2290 fsm_0/nor2_4/a_n37_6# SS0 Vdd Vdd pfet w=6u l=2u
+ ad=12p pd=16u as=0p ps=0u 
M2291 fsm_0/nor2_4/out SA0 fsm_0/nor2_4/a_n37_6# Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2292 fsm_0/nor2_4/out SS0 GND Gnd nfet w=3u l=2u
+ ad=22p pd=20u as=0p ps=0u 
M2293 GND SA0 fsm_0/nor2_4/out Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2294 SA0 fsm_0/inverter_7/in Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2295 SA0 fsm_0/inverter_7/in GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2296 fsm_0/nor2_0/a_n37_6# fsm_0/B2 Vdd Vdd pfet w=6u l=2u
+ ad=12p pd=16u as=0p ps=0u 
M2297 fsm_0/nor2_0/out fsm_0/B1 fsm_0/nor2_0/a_n37_6# Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2298 fsm_0/nor2_0/out fsm_0/B2 GND Gnd nfet w=3u l=2u
+ ad=22p pd=20u as=0p ps=0u 
M2299 GND fsm_0/B1 fsm_0/nor2_0/out Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2300 fsm_0/nor2_2/in2 fsm_0/nor2_0/out Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2301 fsm_0/nor2_2/in2 fsm_0/nor2_0/out GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2302 fsm_0/nor2_1/a_n37_6# fsm_0/B0 Vdd Vdd pfet w=6u l=2u
+ ad=12p pd=16u as=0p ps=0u 
M2303 fsm_0/nor2_1/out fsm_0/B3 fsm_0/nor2_1/a_n37_6# Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2304 fsm_0/nor2_1/out fsm_0/B0 GND Gnd nfet w=3u l=2u
+ ad=22p pd=20u as=0p ps=0u 
M2305 GND fsm_0/B3 fsm_0/nor2_1/out Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2306 fsm_0/nor2_2/in1 fsm_0/nor2_1/out Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2307 fsm_0/nor2_2/in1 fsm_0/nor2_1/out GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2308 fsm_0/nor2_2/a_n37_6# fsm_0/nor2_2/in1 Vdd Vdd pfet w=6u l=2u
+ ad=12p pd=16u as=0p ps=0u 
M2309 fsm_0/nor2_2/out fsm_0/nor2_2/in2 fsm_0/nor2_2/a_n37_6# Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2310 fsm_0/nor2_2/out fsm_0/nor2_2/in1 GND Gnd nfet w=3u l=2u
+ ad=22p pd=20u as=0p ps=0u 
M2311 GND fsm_0/nor2_2/in2 fsm_0/nor2_2/out Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2312 fsm_0/G fsm_0/nor2_2/out Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2313 fsm_0/G fsm_0/nor2_2/out GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2314 fsm_0/nor2_5/a_n37_6# fsm_0/A4 Vdd Vdd pfet w=6u l=2u
+ ad=12p pd=16u as=0p ps=0u 
M2315 fsm_0/nor2_5/out fsm_0/A3 fsm_0/nor2_5/a_n37_6# Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2316 fsm_0/nor2_5/out fsm_0/A4 GND Gnd nfet w=3u l=2u
+ ad=22p pd=20u as=0p ps=0u 
M2317 GND fsm_0/A3 fsm_0/nor2_5/out Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2318 fsm_0/inverter_12/out fsm_0/nor2_5/out Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2319 fsm_0/inverter_12/out fsm_0/nor2_5/out GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2320 fsm_0/inverter_9/in fsm_0/G Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2321 Vdd fsm_0/inverter_12/out fsm_0/inverter_9/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2322 fsm_0/nand2_3/a_n37_n6# fsm_0/G GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2323 fsm_0/inverter_9/in fsm_0/inverter_12/out fsm_0/nand2_3/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2324 fsm_0/inverter_8/in fsm_0/G Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2325 Vdd fsm_0/SR4_0/Q2 fsm_0/inverter_8/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2326 fsm_0/nand2_2/a_n37_n6# fsm_0/G GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2327 fsm_0/inverter_8/in fsm_0/SR4_0/Q2 fsm_0/nand2_2/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2328 fsm_0/inverter_7/in fsm_0/G Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2329 Vdd fsm_0/A1 fsm_0/inverter_7/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2330 fsm_0/nand2_1/a_n37_n6# fsm_0/G GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2331 fsm_0/inverter_7/in fsm_0/A1 fsm_0/nand2_1/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2332 fsm_0/SR4_1/dff3B_2/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2333 fsm_0/SR4_1/dff3B_2/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2334 fsm_0/SR4_1/dff3B_2/gate_0/S fsm_0/SR4_1/dff3B_2/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2335 fsm_0/SR4_1/dff3B_2/gate_0/S fsm_0/SR4_1/dff3B_2/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2336 fsm_0/SR4_1/dff3B_2/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2337 fsm_0/SR4_1/dff3B_2/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2338 fsm_0/SR4_1/dff3B_2/gate_3/Gout fsm_0/B3 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2339 fsm_0/SR4_1/dff3B_2/gate_3/Gout fsm_0/B3 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2340 fsm_0/SR4_1/dff3B_2/gate_3/Gout fsm_0/CLK fsm_0/SR4_1/dff3B_2/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2341 fsm_0/SR4_1/dff3B_2/gate_3/Gout fsm_0/SR4_1/dff3B_2/gate_1/S fsm_0/SR4_1/dff3B_2/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2342 fsm_0/SR4_1/dff3B_2/gate_2/Gout fsm_0/SR4_1/dff3B_2/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2343 fsm_0/SR4_1/dff3B_2/gate_2/Gout fsm_0/SR4_1/dff3B_2/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2344 fsm_0/SR4_1/dff3B_2/gate_2/Gout fsm_0/SR4_1/dff3B_2/gate_2/S fsm_0/SR4_1/dff3B_2/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2345 fsm_0/SR4_1/dff3B_2/gate_2/Gout fsm_0/SR4_1/dff3B_2/gate_0/S fsm_0/SR4_1/dff3B_2/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2346 fsm_0/SR4_1/dff3B_2/Qb fsm_0/B3 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2347 fsm_0/SR4_1/dff3B_2/Qb fsm_0/B3 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2348 fsm_0/B3 fsm_0/SR4_1/dff3B_2/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2349 fsm_0/B3 fsm_0/SR4_1/dff3B_2/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2350 fsm_0/SR4_1/dff3B_2/gate_3/Gin fsm_0/SR4_1/dff3B_2/gate_1/S fsm_0/SR4_1/dff3B_2/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2351 fsm_0/SR4_1/dff3B_2/gate_3/Gin fsm_0/CLK fsm_0/SR4_1/dff3B_2/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2352 fsm_0/SR4_1/dff3B_2/gate_1/Gin fsm_0/SR4_1/dff3B_2/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2353 fsm_0/SR4_1/dff3B_2/gate_1/Gin fsm_0/SR4_1/dff3B_2/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2354 fsm_0/SR4_1/dff3B_2/gate_2/Gin fsm_0/SR4_1/dff3B_2/gate_0/S fsm_0/SR4_1/dff3B_2/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2355 fsm_0/SR4_1/dff3B_2/gate_2/Gin fsm_0/SR4_1/dff3B_2/gate_2/S fsm_0/SR4_1/dff3B_2/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2356 fsm_0/SR4_1/dff3B_2/gate_0/Gin fsm_0/SR4_1/dff3B_2/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2357 fsm_0/SR4_1/dff3B_2/gate_0/Gin fsm_0/SR4_1/dff3B_2/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2358 fsm_0/SR4_1/dff3B_2/inverter_11/in fsm_0/SR4_1/dff3B_2/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2359 Vdd fsm_0/SR4_1/dff3B_2/D fsm_0/SR4_1/dff3B_2/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2360 fsm_0/SR4_1/dff3B_2/nand2_0/a_n37_n6# fsm_0/SR4_1/dff3B_2/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2361 fsm_0/SR4_1/dff3B_2/inverter_11/in fsm_0/SR4_1/dff3B_2/D fsm_0/SR4_1/dff3B_2/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2362 fsm_0/SR4_1/dff3B_2/inverter_7/out RST Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2363 fsm_0/SR4_1/dff3B_2/inverter_7/out RST GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2364 fsm_0/SR4_1/dff3B_2/D fsm_0/SR4_1/S fsm_0/B3 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M2365 fsm_0/SR4_1/dff3B_2/D fsm_0/SR4_1/mux2x1_3/Smb fsm_0/B3 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M2366 fsm_0/SR4_1/dff3B_2/D fsm_0/SR4_1/mux2x1_3/Smb fsm_0/B2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=124p ps=82u 
M2367 fsm_0/SR4_1/dff3B_2/D fsm_0/SR4_1/S fsm_0/B2 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=75p ps=66u 
M2368 fsm_0/SR4_1/mux2x1_3/Smb fsm_0/SR4_1/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2369 fsm_0/SR4_1/mux2x1_3/Smb fsm_0/SR4_1/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2370 fsm_0/SR4_1/dff3B_1/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2371 fsm_0/SR4_1/dff3B_1/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2372 fsm_0/SR4_1/dff3B_1/gate_0/S fsm_0/SR4_1/dff3B_1/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2373 fsm_0/SR4_1/dff3B_1/gate_0/S fsm_0/SR4_1/dff3B_1/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2374 fsm_0/SR4_1/dff3B_1/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2375 fsm_0/SR4_1/dff3B_1/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2376 fsm_0/SR4_1/dff3B_1/gate_3/Gout fsm_0/B2 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2377 fsm_0/SR4_1/dff3B_1/gate_3/Gout fsm_0/B2 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2378 fsm_0/SR4_1/dff3B_1/gate_3/Gout fsm_0/CLK fsm_0/SR4_1/dff3B_1/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2379 fsm_0/SR4_1/dff3B_1/gate_3/Gout fsm_0/SR4_1/dff3B_1/gate_1/S fsm_0/SR4_1/dff3B_1/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2380 fsm_0/SR4_1/dff3B_1/gate_2/Gout fsm_0/SR4_1/dff3B_1/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2381 fsm_0/SR4_1/dff3B_1/gate_2/Gout fsm_0/SR4_1/dff3B_1/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2382 fsm_0/SR4_1/dff3B_1/gate_2/Gout fsm_0/SR4_1/dff3B_1/gate_2/S fsm_0/SR4_1/dff3B_1/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2383 fsm_0/SR4_1/dff3B_1/gate_2/Gout fsm_0/SR4_1/dff3B_1/gate_0/S fsm_0/SR4_1/dff3B_1/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2384 fsm_0/SR4_1/dff3B_1/Qb fsm_0/B2 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2385 fsm_0/SR4_1/dff3B_1/Qb fsm_0/B2 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2386 fsm_0/B2 fsm_0/SR4_1/dff3B_1/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2387 fsm_0/B2 fsm_0/SR4_1/dff3B_1/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2388 fsm_0/SR4_1/dff3B_1/gate_3/Gin fsm_0/SR4_1/dff3B_1/gate_1/S fsm_0/SR4_1/dff3B_1/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2389 fsm_0/SR4_1/dff3B_1/gate_3/Gin fsm_0/CLK fsm_0/SR4_1/dff3B_1/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2390 fsm_0/SR4_1/dff3B_1/gate_1/Gin fsm_0/SR4_1/dff3B_1/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2391 fsm_0/SR4_1/dff3B_1/gate_1/Gin fsm_0/SR4_1/dff3B_1/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2392 fsm_0/SR4_1/dff3B_1/gate_2/Gin fsm_0/SR4_1/dff3B_1/gate_0/S fsm_0/SR4_1/dff3B_1/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2393 fsm_0/SR4_1/dff3B_1/gate_2/Gin fsm_0/SR4_1/dff3B_1/gate_2/S fsm_0/SR4_1/dff3B_1/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2394 fsm_0/SR4_1/dff3B_1/gate_0/Gin fsm_0/SR4_1/dff3B_1/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2395 fsm_0/SR4_1/dff3B_1/gate_0/Gin fsm_0/SR4_1/dff3B_1/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2396 fsm_0/SR4_1/dff3B_1/inverter_11/in fsm_0/SR4_1/dff3B_1/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2397 Vdd fsm_0/SR4_1/dff3B_1/D fsm_0/SR4_1/dff3B_1/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2398 fsm_0/SR4_1/dff3B_1/nand2_0/a_n37_n6# fsm_0/SR4_1/dff3B_1/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2399 fsm_0/SR4_1/dff3B_1/inverter_11/in fsm_0/SR4_1/dff3B_1/D fsm_0/SR4_1/dff3B_1/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2400 fsm_0/SR4_1/dff3B_1/inverter_7/out RST Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2401 fsm_0/SR4_1/dff3B_1/inverter_7/out RST GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2402 fsm_0/SR4_1/dff3B_1/D fsm_0/SR4_1/S fsm_0/B2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M2403 fsm_0/SR4_1/dff3B_1/D fsm_0/SR4_1/mux2x1_2/Smb fsm_0/B2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M2404 fsm_0/SR4_1/dff3B_1/D fsm_0/SR4_1/mux2x1_2/Smb fsm_0/B1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=124p ps=82u 
M2405 fsm_0/SR4_1/dff3B_1/D fsm_0/SR4_1/S fsm_0/B1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=75p ps=66u 
M2406 fsm_0/SR4_1/mux2x1_2/Smb fsm_0/SR4_1/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2407 fsm_0/SR4_1/mux2x1_2/Smb fsm_0/SR4_1/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2408 fsm_0/SR4_1/dff3B_0/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2409 fsm_0/SR4_1/dff3B_0/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2410 fsm_0/SR4_1/dff3B_0/gate_0/S fsm_0/SR4_1/dff3B_0/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2411 fsm_0/SR4_1/dff3B_0/gate_0/S fsm_0/SR4_1/dff3B_0/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2412 fsm_0/SR4_1/dff3B_0/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2413 fsm_0/SR4_1/dff3B_0/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2414 fsm_0/SR4_1/dff3B_0/gate_3/Gout fsm_0/B1 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2415 fsm_0/SR4_1/dff3B_0/gate_3/Gout fsm_0/B1 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2416 fsm_0/SR4_1/dff3B_0/gate_3/Gout fsm_0/CLK fsm_0/SR4_1/dff3B_0/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2417 fsm_0/SR4_1/dff3B_0/gate_3/Gout fsm_0/SR4_1/dff3B_0/gate_1/S fsm_0/SR4_1/dff3B_0/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2418 fsm_0/SR4_1/dff3B_0/gate_2/Gout fsm_0/SR4_1/dff3B_0/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2419 fsm_0/SR4_1/dff3B_0/gate_2/Gout fsm_0/SR4_1/dff3B_0/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2420 fsm_0/SR4_1/dff3B_0/gate_2/Gout fsm_0/SR4_1/dff3B_0/gate_2/S fsm_0/SR4_1/dff3B_0/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2421 fsm_0/SR4_1/dff3B_0/gate_2/Gout fsm_0/SR4_1/dff3B_0/gate_0/S fsm_0/SR4_1/dff3B_0/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2422 fsm_0/SR4_1/dff3B_0/Qb fsm_0/B1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2423 fsm_0/SR4_1/dff3B_0/Qb fsm_0/B1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2424 fsm_0/B1 fsm_0/SR4_1/dff3B_0/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2425 fsm_0/B1 fsm_0/SR4_1/dff3B_0/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2426 fsm_0/SR4_1/dff3B_0/gate_3/Gin fsm_0/SR4_1/dff3B_0/gate_1/S fsm_0/SR4_1/dff3B_0/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2427 fsm_0/SR4_1/dff3B_0/gate_3/Gin fsm_0/CLK fsm_0/SR4_1/dff3B_0/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2428 fsm_0/SR4_1/dff3B_0/gate_1/Gin fsm_0/SR4_1/dff3B_0/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2429 fsm_0/SR4_1/dff3B_0/gate_1/Gin fsm_0/SR4_1/dff3B_0/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2430 fsm_0/SR4_1/dff3B_0/gate_2/Gin fsm_0/SR4_1/dff3B_0/gate_0/S fsm_0/SR4_1/dff3B_0/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2431 fsm_0/SR4_1/dff3B_0/gate_2/Gin fsm_0/SR4_1/dff3B_0/gate_2/S fsm_0/SR4_1/dff3B_0/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2432 fsm_0/SR4_1/dff3B_0/gate_0/Gin fsm_0/SR4_1/dff3B_0/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2433 fsm_0/SR4_1/dff3B_0/gate_0/Gin fsm_0/SR4_1/dff3B_0/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2434 fsm_0/SR4_1/dff3B_0/inverter_11/in fsm_0/SR4_1/dff3B_0/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2435 Vdd fsm_0/SR4_1/dff3B_0/D fsm_0/SR4_1/dff3B_0/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2436 fsm_0/SR4_1/dff3B_0/nand2_0/a_n37_n6# fsm_0/SR4_1/dff3B_0/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2437 fsm_0/SR4_1/dff3B_0/inverter_11/in fsm_0/SR4_1/dff3B_0/D fsm_0/SR4_1/dff3B_0/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2438 fsm_0/SR4_1/dff3B_0/inverter_7/out RST Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2439 fsm_0/SR4_1/dff3B_0/inverter_7/out RST GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2440 fsm_0/SR4_1/dff3B_0/D fsm_0/SR4_1/S fsm_0/B1 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M2441 fsm_0/SR4_1/dff3B_0/D fsm_0/SR4_1/mux2x1_0/Smb fsm_0/B1 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M2442 fsm_0/SR4_1/dff3B_0/D fsm_0/SR4_1/mux2x1_0/Smb fsm_0/B0 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=124p ps=82u 
M2443 fsm_0/SR4_1/dff3B_0/D fsm_0/SR4_1/S fsm_0/B0 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=75p ps=66u 
M2444 fsm_0/SR4_1/dffP_0/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2445 fsm_0/SR4_1/dffP_0/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2446 fsm_0/SR4_1/dffP_0/gate_0/S fsm_0/SR4_1/dffP_0/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2447 fsm_0/SR4_1/dffP_0/gate_0/S fsm_0/SR4_1/dffP_0/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2448 fsm_0/SR4_1/dffP_0/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2449 fsm_0/SR4_1/dffP_0/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2450 fsm_0/SR4_1/dffP_0/gate_3/Gout fsm_0/B0 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2451 fsm_0/SR4_1/dffP_0/gate_3/Gout fsm_0/B0 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2452 fsm_0/SR4_1/dffP_0/gate_3/Gout fsm_0/CLK fsm_0/SR4_1/dffP_0/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2453 fsm_0/SR4_1/dffP_0/gate_3/Gout fsm_0/SR4_1/dffP_0/gate_1/S fsm_0/SR4_1/dffP_0/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2454 fsm_0/SR4_1/dffP_0/gate_2/Gout fsm_0/SR4_1/dffP_0/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2455 fsm_0/SR4_1/dffP_0/gate_2/Gout fsm_0/SR4_1/dffP_0/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2456 fsm_0/SR4_1/dffP_0/gate_2/Gout fsm_0/SR4_1/dffP_0/gate_2/S fsm_0/SR4_1/dffP_0/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2457 fsm_0/SR4_1/dffP_0/gate_2/Gout fsm_0/SR4_1/dffP_0/gate_0/S fsm_0/SR4_1/dffP_0/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2458 fsm_0/SR4_1/dffP_0/Qb fsm_0/B0 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2459 fsm_0/SR4_1/dffP_0/Qb fsm_0/B0 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2460 fsm_0/B0 fsm_0/SR4_1/dffP_0/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2461 fsm_0/B0 fsm_0/SR4_1/dffP_0/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2462 fsm_0/SR4_1/dffP_0/gate_3/Gin fsm_0/SR4_1/dffP_0/gate_1/S fsm_0/SR4_1/dffP_0/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2463 fsm_0/SR4_1/dffP_0/gate_3/Gin fsm_0/CLK fsm_0/SR4_1/dffP_0/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2464 fsm_0/SR4_1/dffP_0/gate_1/Gin fsm_0/SR4_1/dffP_0/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2465 fsm_0/SR4_1/dffP_0/gate_1/Gin fsm_0/SR4_1/dffP_0/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2466 fsm_0/SR4_1/dffP_0/gate_2/Gin fsm_0/SR4_1/dffP_0/gate_0/S fsm_0/SR4_1/dffP_0/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2467 fsm_0/SR4_1/dffP_0/gate_2/Gin fsm_0/SR4_1/dffP_0/gate_2/S fsm_0/SR4_1/dffP_0/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2468 fsm_0/SR4_1/dffP_0/gate_0/Gin fsm_0/SR4_1/dffP_0/nor2_0/out Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2469 fsm_0/SR4_1/dffP_0/gate_0/Gin fsm_0/SR4_1/dffP_0/nor2_0/out GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2470 fsm_0/SR4_1/dffP_0/nor2_0/a_n37_6# RST Vdd Vdd pfet w=6u l=2u
+ ad=12p pd=16u as=0p ps=0u 
M2471 fsm_0/SR4_1/dffP_0/nor2_0/out fsm_0/SR4_1/dffP_0/D fsm_0/SR4_1/dffP_0/nor2_0/a_n37_6# Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2472 fsm_0/SR4_1/dffP_0/nor2_0/out RST GND Gnd nfet w=3u l=2u
+ ad=22p pd=20u as=0p ps=0u 
M2473 GND fsm_0/SR4_1/dffP_0/D fsm_0/SR4_1/dffP_0/nor2_0/out Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2474 fsm_0/SR4_1/dffP_0/D fsm_0/SR4_1/S fsm_0/B0 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M2475 fsm_0/SR4_1/dffP_0/D fsm_0/SR4_1/mux2x1_1/Smb fsm_0/B0 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M2476 fsm_0/SR4_1/dffP_0/D fsm_0/SR4_1/mux2x1_1/Smb fsm_0/SR4_1/INP Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2477 fsm_0/SR4_1/dffP_0/D fsm_0/SR4_1/S fsm_0/SR4_1/INP Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2478 fsm_0/SR4_1/mux2x1_0/Smb fsm_0/SR4_1/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2479 fsm_0/SR4_1/mux2x1_0/Smb fsm_0/SR4_1/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2480 fsm_0/SR4_1/mux2x1_1/Smb fsm_0/SR4_1/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2481 fsm_0/SR4_1/mux2x1_1/Smb fsm_0/SR4_1/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2482 fsm_0/SR4_1/INP fsm_0/B3 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2483 fsm_0/SR4_1/INP fsm_0/B3 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2484 fsm_0/dff3B_0/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2485 fsm_0/dff3B_0/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2486 fsm_0/dff3B_0/gate_0/S fsm_0/dff3B_0/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2487 fsm_0/dff3B_0/gate_0/S fsm_0/dff3B_0/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2488 fsm_0/dff3B_0/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2489 fsm_0/dff3B_0/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2490 fsm_0/dff3B_0/gate_3/Gout fsm_0/A4 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2491 fsm_0/dff3B_0/gate_3/Gout fsm_0/A4 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2492 fsm_0/dff3B_0/gate_3/Gout fsm_0/CLK fsm_0/dff3B_0/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2493 fsm_0/dff3B_0/gate_3/Gout fsm_0/dff3B_0/gate_1/S fsm_0/dff3B_0/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2494 fsm_0/dff3B_0/gate_2/Gout fsm_0/dff3B_0/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2495 fsm_0/dff3B_0/gate_2/Gout fsm_0/dff3B_0/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2496 fsm_0/dff3B_0/gate_2/Gout fsm_0/dff3B_0/gate_2/S fsm_0/dff3B_0/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2497 fsm_0/dff3B_0/gate_2/Gout fsm_0/dff3B_0/gate_0/S fsm_0/dff3B_0/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2498 fsm_0/dff3B_0/Qb fsm_0/A4 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2499 fsm_0/dff3B_0/Qb fsm_0/A4 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2500 fsm_0/A4 fsm_0/dff3B_0/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2501 fsm_0/A4 fsm_0/dff3B_0/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2502 fsm_0/dff3B_0/gate_3/Gin fsm_0/dff3B_0/gate_1/S fsm_0/dff3B_0/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2503 fsm_0/dff3B_0/gate_3/Gin fsm_0/CLK fsm_0/dff3B_0/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2504 fsm_0/dff3B_0/gate_1/Gin fsm_0/dff3B_0/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2505 fsm_0/dff3B_0/gate_1/Gin fsm_0/dff3B_0/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2506 fsm_0/dff3B_0/gate_2/Gin fsm_0/dff3B_0/gate_0/S fsm_0/dff3B_0/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2507 fsm_0/dff3B_0/gate_2/Gin fsm_0/dff3B_0/gate_2/S fsm_0/dff3B_0/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2508 fsm_0/dff3B_0/gate_0/Gin fsm_0/dff3B_0/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2509 fsm_0/dff3B_0/gate_0/Gin fsm_0/dff3B_0/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2510 fsm_0/dff3B_0/inverter_11/in fsm_0/dff3B_0/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2511 Vdd fsm_0/dff3B_0/D fsm_0/dff3B_0/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2512 fsm_0/dff3B_0/nand2_0/a_n37_n6# fsm_0/dff3B_0/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2513 fsm_0/dff3B_0/inverter_11/in fsm_0/dff3B_0/D fsm_0/dff3B_0/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2514 fsm_0/dff3B_0/inverter_7/out RST Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2515 fsm_0/dff3B_0/inverter_7/out RST GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2516 fsm_0/SR4_1/S fsm_0/inverter_2/in Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2517 fsm_0/SR4_1/S fsm_0/inverter_2/in GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2518 fsm_0/inverter_2/in fsm_0/A4 Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2519 Vdd fsm_0/G fsm_0/inverter_2/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2520 fsm_0/nand2_0/a_n37_n6# fsm_0/A4 GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2521 fsm_0/inverter_2/in fsm_0/G fsm_0/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2522 fsm_0/dff3B_0/D fsm_0/SR4_0/S fsm_0/A4 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M2523 fsm_0/dff3B_0/D fsm_0/mux2x1_0/Smb fsm_0/A4 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M2524 fsm_0/dff3B_0/D fsm_0/mux2x1_0/Smb fsm_0/A3 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=124p ps=82u 
M2525 fsm_0/dff3B_0/D fsm_0/SR4_0/S fsm_0/A3 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=75p ps=66u 
M2526 fsm_0/SR4_0/S fsm_0/A4 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2527 fsm_0/SR4_0/S fsm_0/A4 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2528 fsm_0/mux2x1_0/Smb fsm_0/SR4_0/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2529 fsm_0/mux2x1_0/Smb fsm_0/SR4_0/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2530 fsm_0/SR4_0/dff3B_2/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2531 fsm_0/SR4_0/dff3B_2/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2532 fsm_0/SR4_0/dff3B_2/gate_0/S fsm_0/SR4_0/dff3B_2/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2533 fsm_0/SR4_0/dff3B_2/gate_0/S fsm_0/SR4_0/dff3B_2/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2534 fsm_0/SR4_0/dff3B_2/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2535 fsm_0/SR4_0/dff3B_2/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2536 fsm_0/SR4_0/dff3B_2/gate_3/Gout fsm_0/A3 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2537 fsm_0/SR4_0/dff3B_2/gate_3/Gout fsm_0/A3 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2538 fsm_0/SR4_0/dff3B_2/gate_3/Gout fsm_0/CLK fsm_0/SR4_0/dff3B_2/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2539 fsm_0/SR4_0/dff3B_2/gate_3/Gout fsm_0/SR4_0/dff3B_2/gate_1/S fsm_0/SR4_0/dff3B_2/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2540 fsm_0/SR4_0/dff3B_2/gate_2/Gout fsm_0/SR4_0/dff3B_2/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2541 fsm_0/SR4_0/dff3B_2/gate_2/Gout fsm_0/SR4_0/dff3B_2/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2542 fsm_0/SR4_0/dff3B_2/gate_2/Gout fsm_0/SR4_0/dff3B_2/gate_2/S fsm_0/SR4_0/dff3B_2/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2543 fsm_0/SR4_0/dff3B_2/gate_2/Gout fsm_0/SR4_0/dff3B_2/gate_0/S fsm_0/SR4_0/dff3B_2/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2544 fsm_0/SR4_0/dff3B_2/Qb fsm_0/A3 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2545 fsm_0/SR4_0/dff3B_2/Qb fsm_0/A3 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2546 fsm_0/A3 fsm_0/SR4_0/dff3B_2/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2547 fsm_0/A3 fsm_0/SR4_0/dff3B_2/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2548 fsm_0/SR4_0/dff3B_2/gate_3/Gin fsm_0/SR4_0/dff3B_2/gate_1/S fsm_0/SR4_0/dff3B_2/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2549 fsm_0/SR4_0/dff3B_2/gate_3/Gin fsm_0/CLK fsm_0/SR4_0/dff3B_2/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2550 fsm_0/SR4_0/dff3B_2/gate_1/Gin fsm_0/SR4_0/dff3B_2/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2551 fsm_0/SR4_0/dff3B_2/gate_1/Gin fsm_0/SR4_0/dff3B_2/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2552 fsm_0/SR4_0/dff3B_2/gate_2/Gin fsm_0/SR4_0/dff3B_2/gate_0/S fsm_0/SR4_0/dff3B_2/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2553 fsm_0/SR4_0/dff3B_2/gate_2/Gin fsm_0/SR4_0/dff3B_2/gate_2/S fsm_0/SR4_0/dff3B_2/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2554 fsm_0/SR4_0/dff3B_2/gate_0/Gin fsm_0/SR4_0/dff3B_2/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2555 fsm_0/SR4_0/dff3B_2/gate_0/Gin fsm_0/SR4_0/dff3B_2/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2556 fsm_0/SR4_0/dff3B_2/inverter_11/in fsm_0/SR4_0/dff3B_2/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2557 Vdd fsm_0/SR4_0/dff3B_2/D fsm_0/SR4_0/dff3B_2/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2558 fsm_0/SR4_0/dff3B_2/nand2_0/a_n37_n6# fsm_0/SR4_0/dff3B_2/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2559 fsm_0/SR4_0/dff3B_2/inverter_11/in fsm_0/SR4_0/dff3B_2/D fsm_0/SR4_0/dff3B_2/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2560 fsm_0/SR4_0/dff3B_2/inverter_7/out RST Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2561 fsm_0/SR4_0/dff3B_2/inverter_7/out RST GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2562 fsm_0/SR4_0/dff3B_2/D fsm_0/SR4_0/S fsm_0/A3 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M2563 fsm_0/SR4_0/dff3B_2/D fsm_0/SR4_0/mux2x1_3/Smb fsm_0/A3 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M2564 fsm_0/SR4_0/dff3B_2/D fsm_0/SR4_0/mux2x1_3/Smb fsm_0/SR4_0/Q2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=124p ps=82u 
M2565 fsm_0/SR4_0/dff3B_2/D fsm_0/SR4_0/S fsm_0/SR4_0/Q2 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=75p ps=66u 
M2566 fsm_0/SR4_0/mux2x1_3/Smb fsm_0/SR4_0/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2567 fsm_0/SR4_0/mux2x1_3/Smb fsm_0/SR4_0/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2568 fsm_0/SR4_0/dff3B_1/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2569 fsm_0/SR4_0/dff3B_1/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2570 fsm_0/SR4_0/dff3B_1/gate_0/S fsm_0/SR4_0/dff3B_1/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2571 fsm_0/SR4_0/dff3B_1/gate_0/S fsm_0/SR4_0/dff3B_1/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2572 fsm_0/SR4_0/dff3B_1/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2573 fsm_0/SR4_0/dff3B_1/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2574 fsm_0/SR4_0/dff3B_1/gate_3/Gout fsm_0/SR4_0/Q2 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2575 fsm_0/SR4_0/dff3B_1/gate_3/Gout fsm_0/SR4_0/Q2 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2576 fsm_0/SR4_0/dff3B_1/gate_3/Gout fsm_0/CLK fsm_0/SR4_0/dff3B_1/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2577 fsm_0/SR4_0/dff3B_1/gate_3/Gout fsm_0/SR4_0/dff3B_1/gate_1/S fsm_0/SR4_0/dff3B_1/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2578 fsm_0/SR4_0/dff3B_1/gate_2/Gout fsm_0/SR4_0/dff3B_1/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2579 fsm_0/SR4_0/dff3B_1/gate_2/Gout fsm_0/SR4_0/dff3B_1/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2580 fsm_0/SR4_0/dff3B_1/gate_2/Gout fsm_0/SR4_0/dff3B_1/gate_2/S fsm_0/SR4_0/dff3B_1/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2581 fsm_0/SR4_0/dff3B_1/gate_2/Gout fsm_0/SR4_0/dff3B_1/gate_0/S fsm_0/SR4_0/dff3B_1/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2582 fsm_0/SR4_0/dff3B_1/Qb fsm_0/SR4_0/Q2 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2583 fsm_0/SR4_0/dff3B_1/Qb fsm_0/SR4_0/Q2 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2584 fsm_0/SR4_0/Q2 fsm_0/SR4_0/dff3B_1/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2585 fsm_0/SR4_0/Q2 fsm_0/SR4_0/dff3B_1/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2586 fsm_0/SR4_0/dff3B_1/gate_3/Gin fsm_0/SR4_0/dff3B_1/gate_1/S fsm_0/SR4_0/dff3B_1/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2587 fsm_0/SR4_0/dff3B_1/gate_3/Gin fsm_0/CLK fsm_0/SR4_0/dff3B_1/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2588 fsm_0/SR4_0/dff3B_1/gate_1/Gin fsm_0/SR4_0/dff3B_1/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2589 fsm_0/SR4_0/dff3B_1/gate_1/Gin fsm_0/SR4_0/dff3B_1/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2590 fsm_0/SR4_0/dff3B_1/gate_2/Gin fsm_0/SR4_0/dff3B_1/gate_0/S fsm_0/SR4_0/dff3B_1/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2591 fsm_0/SR4_0/dff3B_1/gate_2/Gin fsm_0/SR4_0/dff3B_1/gate_2/S fsm_0/SR4_0/dff3B_1/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2592 fsm_0/SR4_0/dff3B_1/gate_0/Gin fsm_0/SR4_0/dff3B_1/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2593 fsm_0/SR4_0/dff3B_1/gate_0/Gin fsm_0/SR4_0/dff3B_1/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2594 fsm_0/SR4_0/dff3B_1/inverter_11/in fsm_0/SR4_0/dff3B_1/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2595 Vdd fsm_0/SR4_0/dff3B_1/D fsm_0/SR4_0/dff3B_1/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2596 fsm_0/SR4_0/dff3B_1/nand2_0/a_n37_n6# fsm_0/SR4_0/dff3B_1/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2597 fsm_0/SR4_0/dff3B_1/inverter_11/in fsm_0/SR4_0/dff3B_1/D fsm_0/SR4_0/dff3B_1/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2598 fsm_0/SR4_0/dff3B_1/inverter_7/out RST Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2599 fsm_0/SR4_0/dff3B_1/inverter_7/out RST GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2600 fsm_0/SR4_0/dff3B_1/D fsm_0/SR4_0/S fsm_0/SR4_0/Q2 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M2601 fsm_0/SR4_0/dff3B_1/D fsm_0/SR4_0/mux2x1_2/Smb fsm_0/SR4_0/Q2 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M2602 fsm_0/SR4_0/dff3B_1/D fsm_0/SR4_0/mux2x1_2/Smb fsm_0/A1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=124p ps=82u 
M2603 fsm_0/SR4_0/dff3B_1/D fsm_0/SR4_0/S fsm_0/A1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=75p ps=66u 
M2604 fsm_0/SR4_0/mux2x1_2/Smb fsm_0/SR4_0/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2605 fsm_0/SR4_0/mux2x1_2/Smb fsm_0/SR4_0/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2606 fsm_0/SR4_0/dff3B_0/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2607 fsm_0/SR4_0/dff3B_0/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2608 fsm_0/SR4_0/dff3B_0/gate_0/S fsm_0/SR4_0/dff3B_0/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2609 fsm_0/SR4_0/dff3B_0/gate_0/S fsm_0/SR4_0/dff3B_0/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2610 fsm_0/SR4_0/dff3B_0/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2611 fsm_0/SR4_0/dff3B_0/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2612 fsm_0/SR4_0/dff3B_0/gate_3/Gout fsm_0/A1 Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2613 fsm_0/SR4_0/dff3B_0/gate_3/Gout fsm_0/A1 GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2614 fsm_0/SR4_0/dff3B_0/gate_3/Gout fsm_0/CLK fsm_0/SR4_0/dff3B_0/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2615 fsm_0/SR4_0/dff3B_0/gate_3/Gout fsm_0/SR4_0/dff3B_0/gate_1/S fsm_0/SR4_0/dff3B_0/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2616 fsm_0/SR4_0/dff3B_0/gate_2/Gout fsm_0/SR4_0/dff3B_0/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2617 fsm_0/SR4_0/dff3B_0/gate_2/Gout fsm_0/SR4_0/dff3B_0/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2618 fsm_0/SR4_0/dff3B_0/gate_2/Gout fsm_0/SR4_0/dff3B_0/gate_2/S fsm_0/SR4_0/dff3B_0/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2619 fsm_0/SR4_0/dff3B_0/gate_2/Gout fsm_0/SR4_0/dff3B_0/gate_0/S fsm_0/SR4_0/dff3B_0/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2620 fsm_0/SR4_0/dff3B_0/Qb fsm_0/A1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2621 fsm_0/SR4_0/dff3B_0/Qb fsm_0/A1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2622 fsm_0/A1 fsm_0/SR4_0/dff3B_0/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2623 fsm_0/A1 fsm_0/SR4_0/dff3B_0/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2624 fsm_0/SR4_0/dff3B_0/gate_3/Gin fsm_0/SR4_0/dff3B_0/gate_1/S fsm_0/SR4_0/dff3B_0/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2625 fsm_0/SR4_0/dff3B_0/gate_3/Gin fsm_0/CLK fsm_0/SR4_0/dff3B_0/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2626 fsm_0/SR4_0/dff3B_0/gate_1/Gin fsm_0/SR4_0/dff3B_0/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2627 fsm_0/SR4_0/dff3B_0/gate_1/Gin fsm_0/SR4_0/dff3B_0/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2628 fsm_0/SR4_0/dff3B_0/gate_2/Gin fsm_0/SR4_0/dff3B_0/gate_0/S fsm_0/SR4_0/dff3B_0/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2629 fsm_0/SR4_0/dff3B_0/gate_2/Gin fsm_0/SR4_0/dff3B_0/gate_2/S fsm_0/SR4_0/dff3B_0/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2630 fsm_0/SR4_0/dff3B_0/gate_0/Gin fsm_0/SR4_0/dff3B_0/inverter_11/in Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2631 fsm_0/SR4_0/dff3B_0/gate_0/Gin fsm_0/SR4_0/dff3B_0/inverter_11/in GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2632 fsm_0/SR4_0/dff3B_0/inverter_11/in fsm_0/SR4_0/dff3B_0/inverter_7/out Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2633 Vdd fsm_0/SR4_0/dff3B_0/D fsm_0/SR4_0/dff3B_0/inverter_11/in Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2634 fsm_0/SR4_0/dff3B_0/nand2_0/a_n37_n6# fsm_0/SR4_0/dff3B_0/inverter_7/out GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2635 fsm_0/SR4_0/dff3B_0/inverter_11/in fsm_0/SR4_0/dff3B_0/D fsm_0/SR4_0/dff3B_0/nand2_0/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2636 fsm_0/SR4_0/dff3B_0/inverter_7/out RST Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2637 fsm_0/SR4_0/dff3B_0/inverter_7/out RST GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2638 fsm_0/SR4_0/dff3B_0/D fsm_0/SR4_0/S fsm_0/A1 Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M2639 fsm_0/SR4_0/dff3B_0/D fsm_0/SR4_0/mux2x1_0/Smb fsm_0/A1 Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M2640 fsm_0/SR4_0/dff3B_0/D fsm_0/SR4_0/mux2x1_0/Smb fsm_0/CLR Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=124p ps=82u 
M2641 fsm_0/SR4_0/dff3B_0/D fsm_0/SR4_0/S fsm_0/CLR Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=75p ps=66u 
M2642 fsm_0/SR4_0/dffP_0/gate_1/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2643 fsm_0/SR4_0/dffP_0/gate_1/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2644 fsm_0/SR4_0/dffP_0/gate_0/S fsm_0/SR4_0/dffP_0/gate_2/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2645 fsm_0/SR4_0/dffP_0/gate_0/S fsm_0/SR4_0/dffP_0/gate_2/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2646 fsm_0/SR4_0/dffP_0/gate_2/S fsm_0/CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2647 fsm_0/SR4_0/dffP_0/gate_2/S fsm_0/CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2648 fsm_0/SR4_0/dffP_0/gate_3/Gout fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2649 fsm_0/SR4_0/dffP_0/gate_3/Gout fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2650 fsm_0/SR4_0/dffP_0/gate_3/Gout fsm_0/CLK fsm_0/SR4_0/dffP_0/gate_3/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2651 fsm_0/SR4_0/dffP_0/gate_3/Gout fsm_0/SR4_0/dffP_0/gate_1/S fsm_0/SR4_0/dffP_0/gate_3/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2652 fsm_0/SR4_0/dffP_0/gate_2/Gout fsm_0/SR4_0/dffP_0/gate_1/Gin Vdd Vdd pfet w=6u l=2u
+ ad=75p pd=52u as=0p ps=0u 
M2653 fsm_0/SR4_0/dffP_0/gate_2/Gout fsm_0/SR4_0/dffP_0/gate_1/Gin GND Gnd nfet w=3u l=2u
+ ad=47p pd=42u as=0p ps=0u 
M2654 fsm_0/SR4_0/dffP_0/gate_2/Gout fsm_0/SR4_0/dffP_0/gate_2/S fsm_0/SR4_0/dffP_0/gate_2/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=98p ps=60u 
M2655 fsm_0/SR4_0/dffP_0/gate_2/Gout fsm_0/SR4_0/dffP_0/gate_0/S fsm_0/SR4_0/dffP_0/gate_2/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=56p ps=48u 
M2656 fsm_0/SR4_0/dffP_0/Qb fsm_0/CLR Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2657 fsm_0/SR4_0/dffP_0/Qb fsm_0/CLR GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2658 fsm_0/CLR fsm_0/SR4_0/dffP_0/gate_3/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2659 fsm_0/CLR fsm_0/SR4_0/dffP_0/gate_3/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2660 fsm_0/SR4_0/dffP_0/gate_3/Gin fsm_0/SR4_0/dffP_0/gate_1/S fsm_0/SR4_0/dffP_0/gate_1/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2661 fsm_0/SR4_0/dffP_0/gate_3/Gin fsm_0/CLK fsm_0/SR4_0/dffP_0/gate_1/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2662 fsm_0/SR4_0/dffP_0/gate_1/Gin fsm_0/SR4_0/dffP_0/gate_2/Gin Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2663 fsm_0/SR4_0/dffP_0/gate_1/Gin fsm_0/SR4_0/dffP_0/gate_2/Gin GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2664 fsm_0/SR4_0/dffP_0/gate_2/Gin fsm_0/SR4_0/dffP_0/gate_0/S fsm_0/SR4_0/dffP_0/gate_0/Gin Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=75p ps=52u 
M2665 fsm_0/SR4_0/dffP_0/gate_2/Gin fsm_0/SR4_0/dffP_0/gate_2/S fsm_0/SR4_0/dffP_0/gate_0/Gin Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2666 fsm_0/SR4_0/dffP_0/gate_0/Gin fsm_0/SR4_0/dffP_0/nor2_0/out Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2667 fsm_0/SR4_0/dffP_0/gate_0/Gin fsm_0/SR4_0/dffP_0/nor2_0/out GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2668 fsm_0/SR4_0/dffP_0/nor2_0/a_n37_6# RST Vdd Vdd pfet w=6u l=2u
+ ad=12p pd=16u as=0p ps=0u 
M2669 fsm_0/SR4_0/dffP_0/nor2_0/out fsm_0/SR4_0/dffP_0/D fsm_0/SR4_0/dffP_0/nor2_0/a_n37_6# Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2670 fsm_0/SR4_0/dffP_0/nor2_0/out RST GND Gnd nfet w=3u l=2u
+ ad=22p pd=20u as=0p ps=0u 
M2671 GND fsm_0/SR4_0/dffP_0/D fsm_0/SR4_0/dffP_0/nor2_0/out Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2672 fsm_0/SR4_0/dffP_0/D fsm_0/SR4_0/S fsm_0/CLR Vdd pfet w=6u l=2u
+ ad=98p pd=60u as=0p ps=0u 
M2673 fsm_0/SR4_0/dffP_0/D fsm_0/SR4_0/mux2x1_1/Smb fsm_0/CLR Gnd nfet w=3u l=2u
+ ad=56p pd=48u as=0p ps=0u 
M2674 fsm_0/SR4_0/dffP_0/D fsm_0/SR4_0/mux2x1_1/Smb fsm_0/SS1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=85p ps=54u 
M2675 fsm_0/SR4_0/dffP_0/D fsm_0/SR4_0/S fsm_0/SS1 Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=47p ps=42u 
M2676 fsm_0/SR4_0/mux2x1_0/Smb fsm_0/SR4_0/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2677 fsm_0/SR4_0/mux2x1_0/Smb fsm_0/SR4_0/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2678 fsm_0/SR4_0/mux2x1_1/Smb fsm_0/SR4_0/S Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2679 fsm_0/SR4_0/mux2x1_1/Smb fsm_0/SR4_0/S GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2680 fsm_0/SS1 fsm_0/xor2_0/nand2_4/nand_in1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2681 Vdd fsm_0/xor2_0/nand2_4/nand_in2 fsm_0/SS1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2682 fsm_0/xor2_0/nand2_4/a_n37_n6# fsm_0/xor2_0/nand2_4/nand_in1 GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2683 fsm_0/SS1 fsm_0/xor2_0/nand2_4/nand_in2 fsm_0/xor2_0/nand2_4/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2684 fsm_0/xor2_0/nand2_4/nand_in1 fsm_0/SR4_0/S Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2685 Vdd fsm_0/xor2_0/nand2_3/nand_in2 fsm_0/xor2_0/nand2_4/nand_in1 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2686 fsm_0/xor2_0/nand2_3/a_n37_n6# fsm_0/SR4_0/S GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2687 fsm_0/xor2_0/nand2_4/nand_in1 fsm_0/xor2_0/nand2_3/nand_in2 fsm_0/xor2_0/nand2_3/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2688 fsm_0/xor2_0/nand2_4/nand_in2 fsm_0/xor2_0/nand2_3/nand_in2 Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2689 Vdd fsm_0/SR4_0/S fsm_0/xor2_0/nand2_4/nand_in2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2690 fsm_0/xor2_0/nand2_2/a_n37_n6# fsm_0/xor2_0/nand2_3/nand_in2 GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2691 fsm_0/xor2_0/nand2_4/nand_in2 fsm_0/SR4_0/S fsm_0/xor2_0/nand2_2/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2692 fsm_0/xor2_0/nand2_3/nand_in2 fsm_0/SR4_0/S Vdd Vdd pfet w=6u l=2u
+ ad=36p pd=24u as=0p ps=0u 
M2693 Vdd fsm_0/SR4_0/S fsm_0/xor2_0/nand2_3/nand_in2 Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M2694 fsm_0/xor2_0/nand2_1/a_n37_n6# fsm_0/SR4_0/S GND Gnd nfet w=3u l=2u
+ ad=6p pd=10u as=0p ps=0u 
M2695 fsm_0/xor2_0/nand2_3/nand_in2 fsm_0/SR4_0/S fsm_0/xor2_0/nand2_1/a_n37_n6# Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2696 fsm_0/CLK inverter_1/in Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2697 fsm_0/CLK inverter_1/in GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
M2698 inverter_1/in CLK Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=0p ps=0u 
M2699 inverter_1/in CLK GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=0p ps=0u 
C0 SA0 Vdd 2.3fF
C1 Vdd fsm_0/A3 6.3fF
C2 Vdd fsm_0/A1 5.0fF
C3 Vdd fsm_0/CLK 33.4fF
C4 Vdd SB0 2.3fF
C5 Vdd fsm_0/B1 5.3fF
C6 SA0 SA1 3.1fF
C7 Vdd SB1 2.6fF
C8 fsm_0/SR4_0/Q2 Vdd 5.3fF
C9 Vdd SA1 2.3fF
C10 SS0 fsm_0/CLR 2.2fF
C11 fsm_0/B0 Vdd 2.8fF
C12 nor2_0/in2 Vdd 2.2fF
C13 Vdd fsm_0/B2 5.4fF
C14 fsm_0/CLK fsm_0/CLR 2.8fF
C15 Vdd fsm_0/CLR 16.5fF
C16 Vdd fsm_0/B3 5.8fF
C17 Vdd SS0 6.0fF
C18 SubB_0/QB0 Vdd 2.1fF
C19 CLK gnd! 5.2fF
C20 inverter_1/in gnd! 8.3fF
C21 fsm_0/xor2_0/nand2_3/nand_in2 gnd! 28.1fF
C22 fsm_0/xor2_0/nand2_4/nand_in2 gnd! 17.8fF
C23 fsm_0/xor2_0/nand2_4/nand_in1 gnd! 12.2fF
C24 fsm_0/SS1 gnd! 9.9fF
C25 fsm_0/SR4_0/mux2x1_1/Smb gnd! 20.4fF
C26 fsm_0/SR4_0/dffP_0/D gnd! 13.4fF
C27 fsm_0/SR4_0/dffP_0/nor2_0/out gnd! 9.3fF
C28 fsm_0/SR4_0/dffP_0/gate_0/Gin gnd! 6.2fF
C29 fsm_0/SR4_0/dffP_0/Qb gnd! 2.1fF
C30 fsm_0/SR4_0/dffP_0/gate_2/Gin gnd! 16.9fF
C31 fsm_0/SR4_0/dffP_0/gate_2/Gout gnd! 4.4fF
C32 fsm_0/SR4_0/dffP_0/gate_1/Gin gnd! 17.3fF
C33 fsm_0/SR4_0/dffP_0/gate_3/Gin gnd! 17.4fF
C34 fsm_0/SR4_0/dffP_0/gate_3/Gout gnd! 4.4fF
C35 fsm_0/SR4_0/dffP_0/gate_0/S gnd! 26.8fF
C36 fsm_0/SR4_0/dffP_0/gate_2/S gnd! 33.8fF
C37 fsm_0/SR4_0/dffP_0/gate_1/S gnd! 27.0fF
C38 fsm_0/CLR gnd! 708.3fF
C39 fsm_0/SR4_0/mux2x1_0/Smb gnd! 20.4fF
C40 fsm_0/SR4_0/dff3B_0/D gnd! 15.5fF
C41 fsm_0/SR4_0/dff3B_0/inverter_7/out gnd! 11.5fF
C42 fsm_0/SR4_0/dff3B_0/inverter_11/in gnd! 10.5fF
C43 fsm_0/SR4_0/dff3B_0/gate_0/Gin gnd! 6.2fF
C44 fsm_0/SR4_0/dff3B_0/Qb gnd! 2.1fF
C45 fsm_0/SR4_0/dff3B_0/gate_2/Gin gnd! 16.9fF
C46 fsm_0/SR4_0/dff3B_0/gate_2/Gout gnd! 4.4fF
C47 fsm_0/SR4_0/dff3B_0/gate_1/Gin gnd! 17.3fF
C48 fsm_0/SR4_0/dff3B_0/gate_3/Gin gnd! 17.4fF
C49 fsm_0/SR4_0/dff3B_0/gate_3/Gout gnd! 4.4fF
C50 fsm_0/SR4_0/dff3B_0/gate_0/S gnd! 26.8fF
C51 fsm_0/SR4_0/dff3B_0/gate_2/S gnd! 33.8fF
C52 fsm_0/SR4_0/dff3B_0/gate_1/S gnd! 26.8fF
C53 fsm_0/SR4_0/mux2x1_2/Smb gnd! 20.4fF
C54 fsm_0/SR4_0/dff3B_1/D gnd! 15.5fF
C55 fsm_0/SR4_0/dff3B_1/inverter_7/out gnd! 11.5fF
C56 fsm_0/SR4_0/dff3B_1/inverter_11/in gnd! 10.5fF
C57 fsm_0/SR4_0/dff3B_1/gate_0/Gin gnd! 6.2fF
C58 fsm_0/SR4_0/dff3B_1/Qb gnd! 2.1fF
C59 fsm_0/SR4_0/dff3B_1/gate_2/Gin gnd! 16.9fF
C60 fsm_0/SR4_0/dff3B_1/gate_2/Gout gnd! 4.4fF
C61 fsm_0/SR4_0/dff3B_1/gate_1/Gin gnd! 17.3fF
C62 fsm_0/SR4_0/dff3B_1/gate_3/Gin gnd! 17.4fF
C63 fsm_0/SR4_0/dff3B_1/gate_3/Gout gnd! 4.4fF
C64 fsm_0/SR4_0/dff3B_1/gate_0/S gnd! 26.8fF
C65 fsm_0/SR4_0/dff3B_1/gate_2/S gnd! 33.8fF
C66 fsm_0/SR4_0/dff3B_1/gate_1/S gnd! 26.8fF
C67 fsm_0/SR4_0/mux2x1_3/Smb gnd! 20.4fF
C68 fsm_0/SR4_0/dff3B_2/D gnd! 15.5fF
C69 fsm_0/SR4_0/dff3B_2/inverter_7/out gnd! 11.5fF
C70 fsm_0/SR4_0/dff3B_2/inverter_11/in gnd! 10.5fF
C71 fsm_0/SR4_0/dff3B_2/gate_0/Gin gnd! 6.2fF
C72 fsm_0/SR4_0/dff3B_2/Qb gnd! 2.1fF
C73 fsm_0/SR4_0/dff3B_2/gate_2/Gin gnd! 16.9fF
C74 fsm_0/SR4_0/dff3B_2/gate_2/Gout gnd! 4.4fF
C75 fsm_0/SR4_0/dff3B_2/gate_1/Gin gnd! 17.3fF
C76 fsm_0/SR4_0/dff3B_2/gate_3/Gin gnd! 17.4fF
C77 fsm_0/SR4_0/dff3B_2/gate_3/Gout gnd! 4.4fF
C78 fsm_0/SR4_0/dff3B_2/gate_0/S gnd! 26.8fF
C79 fsm_0/SR4_0/dff3B_2/gate_2/S gnd! 33.8fF
C80 fsm_0/SR4_0/dff3B_2/gate_1/S gnd! 26.8fF
C81 fsm_0/SR4_0/S gnd! 256.3fF
C82 fsm_0/A3 gnd! 186.3fF
C83 fsm_0/mux2x1_0/Smb gnd! 20.3fF
C84 fsm_0/G gnd! 87.0fF
C85 fsm_0/A4 gnd! 100.8fF
C86 fsm_0/inverter_2/in gnd! 9.8fF
C87 fsm_0/dff3B_0/D gnd! 15.4fF
C88 fsm_0/dff3B_0/inverter_7/out gnd! 11.5fF
C89 fsm_0/dff3B_0/inverter_11/in gnd! 10.5fF
C90 fsm_0/dff3B_0/gate_0/Gin gnd! 6.2fF
C91 fsm_0/dff3B_0/Qb gnd! 2.1fF
C92 fsm_0/dff3B_0/gate_2/Gin gnd! 16.9fF
C93 fsm_0/dff3B_0/gate_2/Gout gnd! 4.4fF
C94 fsm_0/dff3B_0/gate_1/Gin gnd! 17.3fF
C95 fsm_0/dff3B_0/gate_3/Gin gnd! 17.4fF
C96 fsm_0/dff3B_0/gate_3/Gout gnd! 4.4fF
C97 fsm_0/dff3B_0/gate_0/S gnd! 26.8fF
C98 fsm_0/dff3B_0/gate_2/S gnd! 33.8fF
C99 fsm_0/dff3B_0/gate_1/S gnd! 26.8fF
C100 fsm_0/CLK gnd! 2471.7fF
C101 fsm_0/B3 gnd! 173.1fF
C102 fsm_0/SR4_1/INP gnd! 6.2fF
C103 fsm_0/SR4_1/mux2x1_1/Smb gnd! 20.4fF
C104 fsm_0/SR4_1/dffP_0/D gnd! 13.4fF
C105 fsm_0/SR4_1/dffP_0/nor2_0/out gnd! 9.3fF
C106 fsm_0/SR4_1/dffP_0/gate_0/Gin gnd! 6.2fF
C107 fsm_0/SR4_1/dffP_0/Qb gnd! 2.1fF
C108 fsm_0/SR4_1/dffP_0/gate_2/Gin gnd! 16.9fF
C109 fsm_0/SR4_1/dffP_0/gate_2/Gout gnd! 4.4fF
C110 fsm_0/SR4_1/dffP_0/gate_1/Gin gnd! 17.3fF
C111 fsm_0/SR4_1/dffP_0/gate_3/Gin gnd! 17.4fF
C112 fsm_0/SR4_1/dffP_0/gate_3/Gout gnd! 4.4fF
C113 fsm_0/SR4_1/dffP_0/gate_0/S gnd! 26.8fF
C114 fsm_0/SR4_1/dffP_0/gate_2/S gnd! 33.8fF
C115 fsm_0/SR4_1/dffP_0/gate_1/S gnd! 26.8fF
C116 fsm_0/SR4_1/mux2x1_0/Smb gnd! 20.4fF
C117 fsm_0/SR4_1/dff3B_0/D gnd! 15.5fF
C118 fsm_0/SR4_1/dff3B_0/inverter_7/out gnd! 11.5fF
C119 fsm_0/SR4_1/dff3B_0/inverter_11/in gnd! 10.5fF
C120 fsm_0/SR4_1/dff3B_0/gate_0/Gin gnd! 6.2fF
C121 fsm_0/SR4_1/dff3B_0/Qb gnd! 2.1fF
C122 fsm_0/SR4_1/dff3B_0/gate_2/Gin gnd! 16.9fF
C123 fsm_0/SR4_1/dff3B_0/gate_2/Gout gnd! 4.4fF
C124 fsm_0/SR4_1/dff3B_0/gate_1/Gin gnd! 17.3fF
C125 fsm_0/SR4_1/dff3B_0/gate_3/Gin gnd! 17.4fF
C126 fsm_0/SR4_1/dff3B_0/gate_3/Gout gnd! 4.4fF
C127 fsm_0/SR4_1/dff3B_0/gate_0/S gnd! 26.8fF
C128 fsm_0/SR4_1/dff3B_0/gate_2/S gnd! 33.8fF
C129 fsm_0/SR4_1/dff3B_0/gate_1/S gnd! 27.0fF
C130 fsm_0/B1 gnd! 113.0fF
C131 fsm_0/SR4_1/mux2x1_2/Smb gnd! 20.4fF
C132 fsm_0/SR4_1/dff3B_1/D gnd! 15.5fF
C133 fsm_0/SR4_1/dff3B_1/inverter_7/out gnd! 11.5fF
C134 fsm_0/SR4_1/dff3B_1/inverter_11/in gnd! 10.5fF
C135 fsm_0/SR4_1/dff3B_1/gate_0/Gin gnd! 6.2fF
C136 fsm_0/SR4_1/dff3B_1/Qb gnd! 2.1fF
C137 fsm_0/SR4_1/dff3B_1/gate_2/Gin gnd! 16.9fF
C138 fsm_0/SR4_1/dff3B_1/gate_2/Gout gnd! 4.4fF
C139 fsm_0/SR4_1/dff3B_1/gate_1/Gin gnd! 17.3fF
C140 fsm_0/SR4_1/dff3B_1/gate_3/Gin gnd! 17.4fF
C141 fsm_0/SR4_1/dff3B_1/gate_3/Gout gnd! 4.4fF
C142 fsm_0/SR4_1/dff3B_1/gate_0/S gnd! 26.8fF
C143 fsm_0/SR4_1/dff3B_1/gate_2/S gnd! 33.8fF
C144 fsm_0/SR4_1/dff3B_1/gate_1/S gnd! 26.8fF
C145 fsm_0/B2 gnd! 118.3fF
C146 fsm_0/SR4_1/mux2x1_3/Smb gnd! 20.4fF
C147 fsm_0/SR4_1/S gnd! 156.9fF
C148 RST gnd! 231.9fF
C149 fsm_0/SR4_1/dff3B_2/D gnd! 15.5fF
C150 fsm_0/SR4_1/dff3B_2/inverter_7/out gnd! 11.5fF
C151 fsm_0/SR4_1/dff3B_2/inverter_11/in gnd! 10.5fF
C152 fsm_0/SR4_1/dff3B_2/gate_0/Gin gnd! 6.2fF
C153 fsm_0/SR4_1/dff3B_2/Qb gnd! 2.1fF
C154 fsm_0/SR4_1/dff3B_2/gate_2/Gin gnd! 16.9fF
C155 fsm_0/SR4_1/dff3B_2/gate_2/Gout gnd! 4.4fF
C156 fsm_0/SR4_1/dff3B_2/gate_1/Gin gnd! 17.3fF
C157 fsm_0/SR4_1/dff3B_2/gate_3/Gin gnd! 17.4fF
C158 fsm_0/SR4_1/dff3B_2/gate_3/Gout gnd! 4.4fF
C159 Vdd gnd! 1299.7fF
C160 fsm_0/SR4_1/dff3B_2/gate_0/S gnd! 26.8fF
C161 fsm_0/SR4_1/dff3B_2/gate_2/S gnd! 33.8fF
C162 fsm_0/SR4_1/dff3B_2/gate_1/S gnd! 26.8fF
C163 fsm_0/A1 gnd! 112.4fF
C164 fsm_0/SR4_0/Q2 gnd! 108.3fF
C165 fsm_0/inverter_12/out gnd! 11.0fF
C166 fsm_0/nor2_5/out gnd! 9.5fF
C167 fsm_0/nor2_2/out gnd! 9.2fF
C168 fsm_0/nor2_2/in1 gnd! 8.8fF
C169 fsm_0/nor2_1/out gnd! 9.2fF
C170 fsm_0/B0 gnd! 105.2fF
C171 fsm_0/nor2_2/in2 gnd! 19.2fF
C172 fsm_0/nor2_0/out gnd! 9.2fF
C173 fsm_0/inverter_7/in gnd! 10.4fF
C174 SA0 gnd! 351.6fF
C175 fsm_0/inverter_8/in gnd! 10.4fF
C176 SB0 gnd! 419.9fF
C177 SS0 gnd! 415.7fF
C178 fsm_0/inverter_9/in gnd! 10.4fF
C179 SA1 gnd! 448.8fF
C180 fsm_0/nor2_4/out gnd! 11.0fF
C181 SB1 gnd! 526.3fF
C182 fsm_0/nor2_3/out gnd! 11.0fF
C183 nor2_0/in2 gnd! 35.6fF
C184 nor2_0/in1 gnd! 8.4fF
C185 SubB_0/dff3B_0/Q gnd! 85.7fF
C186 SubB_0/mux2x1_0/Sm gnd! 17.5fF
C187 AbS gnd! 75.4fF
C188 SubB_0/abs_0/xor2_0/nand2_3/nand_in2 gnd! 28.1fF
C189 SubB_0/abs_0/xor2_0/nand2_4/nand_in2 gnd! 17.8fF
C190 SubB_0/abs_0/xor2_0/nand2_4/nand_in1 gnd! 12.2fF
C191 SubB_0/abs_0/ha_0/not1_0/not_in gnd! 9.8fF
C192 SubB_0/abs_0/ha_0/ha_in2 gnd! 48.0fF
C193 SubB_0/abs_0/ha_0/xor2_0/nand2_3/nand_in2 gnd! 28.1fF
C194 SubB_0/abs_0/ha_0/xor2_0/nand2_4/nand_in2 gnd! 17.8fF
C195 SubB_0/abs_0/ha_0/xor2_0/nand2_4/nand_in1 gnd! 12.2fF
C196 SubB_0/abs_0/ha_1/not1_0/not_in gnd! 9.8fF
C197 SubB_0/abs_0/cin gnd! 48.0fF
C198 SubB_0/abs_0/ha_1/xor2_0/nand2_3/nand_in2 gnd! 28.1fF
C199 SubB_0/abs_0/ha_1/ha_in1 gnd! 36.9fF
C200 SubB_0/abs_0/sum gnd! 114.7fF
C201 SubB_0/abs_0/ha_1/xor2_0/nand2_4/nand_in2 gnd! 17.8fF
C202 SubB_0/abs_0/ha_1/xor2_0/nand2_4/nand_in1 gnd! 12.2fF
C203 SubB_0/abs_0/nor2_0/in2 gnd! 16.5fF
C204 SubB_0/abs_0/nor2_0/in1 gnd! 21.2fF
C205 SubB_0/dff3B_0/D gnd! 69.3fF
C206 SubB_0/abs_0/nor2_0/out gnd! 8.8fF
C207 SubB_0/SR2B_0/mux4x1_0/mux2x1_1/Smb gnd! 39.1fF
C208 SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Smb gnd! 22.7fF
C209 A0 gnd! 3.7fF
C210 SR gnd! 3.7fF
C211 SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Min1 gnd! 9.7fF
C212 SubB_0/SR2B_0/mux4x1_0/mux2x1_2/Min2 gnd! 12.2fF
C213 SubB_0/SR2B_0/mux4x1_1/mux2x1_1/Smb gnd! 39.5fF
C214 SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Smb gnd! 22.7fF
C215 A1 gnd! 3.7fF
C216 SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Min1 gnd! 9.7fF
C217 SubB_0/SR2B_0/mux4x1_1/mux2x1_2/Min2 gnd! 12.2fF
C218 SubB_0/SR2B_0/mux4x1_2/mux2x1_1/Smb gnd! 39.1fF
C219 SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Smb gnd! 22.7fF
C220 A2 gnd! 3.7fF
C221 SubB_0/SR2B_0/Q1 gnd! 147.3fF
C222 SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Min1 gnd! 9.7fF
C223 SubB_0/SR2B_0/mux4x1_2/mux2x1_2/Min2 gnd! 12.2fF
C224 SubB_0/SR2B_0/mux4x1_3/mux2x1_1/Smb gnd! 39.1fF
C225 SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Smb gnd! 22.7fF
C226 A3 gnd! 3.7fF
C227 SubB_0/SR2B_0/Q2 gnd! 134.6fF
C228 SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Min1 gnd! 9.7fF
C229 SubB_0/SR2B_0/mux4x1_3/mux2x1_2/Min2 gnd! 12.2fF
C230 SubB_0/SR2B_0/mux4x1_4/mux2x1_1/Smb gnd! 39.1fF
C231 SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Smb gnd! 22.7fF
C232 A4 gnd! 3.7fF
C233 SubB_0/SR2B_0/Q3 gnd! 146.9fF
C234 SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Min1 gnd! 9.7fF
C235 SubB_0/SR2B_0/mux4x1_4/mux2x1_2/Min2 gnd! 12.2fF
C236 SubB_0/SR2B_0/mux4x1_5/mux2x1_1/Smb gnd! 39.1fF
C237 SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Smb gnd! 22.7fF
C238 A5 gnd! 3.7fF
C239 SubB_0/SR2B_0/Q4 gnd! 134.6fF
C240 SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Min1 gnd! 9.7fF
C241 SubB_0/SR2B_0/mux4x1_5/mux2x1_2/Min2 gnd! 12.2fF
C242 SubB_0/SR2B_0/mux4x1_6/mux2x1_1/Smb gnd! 39.1fF
C243 SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Smb gnd! 22.7fF
C244 A6 gnd! 3.7fF
C245 SubB_0/SR2B_0/Q5 gnd! 118.7fF
C246 SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Min1 gnd! 9.7fF
C247 SubB_0/SR2B_0/mux4x1_6/mux2x1_2/Min2 gnd! 12.2fF
C248 SubB_0/SR2B_0/mux4x1_7/mux2x1_1/Smb gnd! 39.1fF
C249 SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Smb gnd! 22.7fF
C250 A7 gnd! 3.7fF
C251 SubB_0/SR2B_0/Q6 gnd! 134.6fF
C252 SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Min1 gnd! 9.7fF
C253 SubB_0/QA0 gnd! 249.6fF
C254 SubB_0/SR2B_0/mux4x1_7/mux2x1_2/Min2 gnd! 12.2fF
C255 SubB_0/SR2B_0/Q7 gnd! 115.7fF
C256 SubB_0/SR2B_0/dff3B_0/D gnd! 21.7fF
C257 SubB_0/SR2B_0/dff3B_0/inverter_7/out gnd! 11.5fF
C258 SubB_0/SR2B_0/dff3B_0/inverter_11/in gnd! 10.5fF
C259 SubB_0/SR2B_0/dff3B_0/gate_0/Gin gnd! 6.2fF
C260 SubB_0/SR2B_0/dff3B_0/Qb gnd! 2.1fF
C261 SubB_0/SR2B_0/dff3B_0/gate_2/Gin gnd! 16.9fF
C262 SubB_0/SR2B_0/dff3B_0/gate_2/Gout gnd! 4.4fF
C263 SubB_0/SR2B_0/dff3B_0/gate_1/Gin gnd! 17.3fF
C264 SubB_0/SR2B_0/dff3B_0/gate_3/Gin gnd! 17.4fF
C265 SubB_0/SR2B_0/dff3B_0/gate_3/Gout gnd! 4.4fF
C266 SubB_0/SR2B_0/dff3B_0/gate_0/S gnd! 26.8fF
C267 SubB_0/SR2B_0/dff3B_0/gate_2/S gnd! 33.8fF
C268 SubB_0/SR2B_0/dff3B_0/gate_1/S gnd! 27.4fF
C269 SubB_0/SR2B_0/dff3B_1/D gnd! 21.7fF
C270 SubB_0/SR2B_0/dff3B_1/inverter_7/out gnd! 11.5fF
C271 SubB_0/SR2B_0/dff3B_1/inverter_11/in gnd! 10.5fF
C272 SubB_0/SR2B_0/dff3B_1/gate_0/Gin gnd! 6.2fF
C273 SubB_0/SR2B_0/dff3B_1/Qb gnd! 2.1fF
C274 SubB_0/SR2B_0/dff3B_1/gate_2/Gin gnd! 16.9fF
C275 SubB_0/SR2B_0/dff3B_1/gate_2/Gout gnd! 4.4fF
C276 SubB_0/SR2B_0/dff3B_1/gate_1/Gin gnd! 17.3fF
C277 SubB_0/SR2B_0/dff3B_1/gate_3/Gin gnd! 17.4fF
C278 SubB_0/SR2B_0/dff3B_1/gate_3/Gout gnd! 4.4fF
C279 SubB_0/SR2B_0/dff3B_1/gate_0/S gnd! 26.8fF
C280 SubB_0/SR2B_0/dff3B_1/gate_2/S gnd! 33.8fF
C281 SubB_0/SR2B_0/dff3B_1/gate_1/S gnd! 27.4fF
C282 SubB_0/SR2B_0/dff3B_2/D gnd! 21.7fF
C283 SubB_0/SR2B_0/dff3B_2/inverter_7/out gnd! 11.5fF
C284 SubB_0/SR2B_0/dff3B_2/inverter_11/in gnd! 10.5fF
C285 SubB_0/SR2B_0/dff3B_2/gate_0/Gin gnd! 6.2fF
C286 SubB_0/SR2B_0/dff3B_2/Qb gnd! 2.1fF
C287 SubB_0/SR2B_0/dff3B_2/gate_2/Gin gnd! 16.9fF
C288 SubB_0/SR2B_0/dff3B_2/gate_2/Gout gnd! 4.4fF
C289 SubB_0/SR2B_0/dff3B_2/gate_1/Gin gnd! 17.3fF
C290 SubB_0/SR2B_0/dff3B_2/gate_3/Gin gnd! 17.4fF
C291 SubB_0/SR2B_0/dff3B_2/gate_3/Gout gnd! 4.4fF
C292 SubB_0/SR2B_0/dff3B_2/gate_0/S gnd! 26.8fF
C293 SubB_0/SR2B_0/dff3B_2/gate_2/S gnd! 33.8fF
C294 SubB_0/SR2B_0/dff3B_2/gate_1/S gnd! 27.4fF
C295 SubB_0/SR2B_0/dff3B_3/D gnd! 21.7fF
C296 SubB_0/SR2B_0/dff3B_3/inverter_7/out gnd! 11.5fF
C297 SubB_0/SR2B_0/dff3B_3/inverter_11/in gnd! 10.5fF
C298 SubB_0/SR2B_0/dff3B_3/gate_0/Gin gnd! 6.2fF
C299 SubB_0/SR2B_0/dff3B_3/Qb gnd! 2.1fF
C300 SubB_0/SR2B_0/dff3B_3/gate_2/Gin gnd! 16.9fF
C301 SubB_0/SR2B_0/dff3B_3/gate_2/Gout gnd! 4.4fF
C302 SubB_0/SR2B_0/dff3B_3/gate_1/Gin gnd! 17.3fF
C303 SubB_0/SR2B_0/dff3B_3/gate_3/Gin gnd! 17.4fF
C304 SubB_0/SR2B_0/dff3B_3/gate_3/Gout gnd! 4.4fF
C305 SubB_0/SR2B_0/dff3B_3/gate_0/S gnd! 26.8fF
C306 SubB_0/SR2B_0/dff3B_3/gate_2/S gnd! 33.8fF
C307 SubB_0/SR2B_0/dff3B_3/gate_1/S gnd! 27.4fF
C308 SubB_0/SR2B_0/dff3B_4/D gnd! 21.7fF
C309 SubB_0/SR2B_0/dff3B_4/inverter_7/out gnd! 11.5fF
C310 SubB_0/SR2B_0/dff3B_4/inverter_11/in gnd! 10.5fF
C311 SubB_0/SR2B_0/dff3B_4/gate_0/Gin gnd! 6.2fF
C312 SubB_0/SR2B_0/dff3B_4/Qb gnd! 2.1fF
C313 SubB_0/SR2B_0/dff3B_4/gate_2/Gin gnd! 16.9fF
C314 SubB_0/SR2B_0/dff3B_4/gate_2/Gout gnd! 4.4fF
C315 SubB_0/SR2B_0/dff3B_4/gate_1/Gin gnd! 17.3fF
C316 SubB_0/SR2B_0/dff3B_4/gate_3/Gin gnd! 17.4fF
C317 SubB_0/SR2B_0/dff3B_4/gate_3/Gout gnd! 4.4fF
C318 SubB_0/SR2B_0/dff3B_4/gate_0/S gnd! 26.8fF
C319 SubB_0/SR2B_0/dff3B_4/gate_2/S gnd! 33.8fF
C320 SubB_0/SR2B_0/dff3B_4/gate_1/S gnd! 27.4fF
C321 SubB_0/SR2B_0/dff3B_5/D gnd! 21.7fF
C322 SubB_0/SR2B_0/dff3B_5/inverter_7/out gnd! 11.5fF
C323 SubB_0/SR2B_0/dff3B_5/inverter_11/in gnd! 10.5fF
C324 SubB_0/SR2B_0/dff3B_5/gate_0/Gin gnd! 6.2fF
C325 SubB_0/SR2B_0/dff3B_5/Qb gnd! 2.1fF
C326 SubB_0/SR2B_0/dff3B_5/gate_2/Gin gnd! 16.9fF
C327 SubB_0/SR2B_0/dff3B_5/gate_2/Gout gnd! 4.4fF
C328 SubB_0/SR2B_0/dff3B_5/gate_1/Gin gnd! 17.3fF
C329 SubB_0/SR2B_0/dff3B_5/gate_3/Gin gnd! 17.4fF
C330 SubB_0/SR2B_0/dff3B_5/gate_3/Gout gnd! 4.4fF
C331 SubB_0/SR2B_0/dff3B_5/gate_0/S gnd! 26.8fF
C332 SubB_0/SR2B_0/dff3B_5/gate_2/S gnd! 33.8fF
C333 SubB_0/SR2B_0/dff3B_5/gate_1/S gnd! 27.4fF
C334 SubB_0/SR2B_0/dff3B_6/D gnd! 21.7fF
C335 SubB_0/SR2B_0/dff3B_6/inverter_7/out gnd! 11.5fF
C336 SubB_0/SR2B_0/dff3B_6/inverter_11/in gnd! 10.5fF
C337 SubB_0/SR2B_0/dff3B_6/gate_0/Gin gnd! 6.2fF
C338 SubB_0/SR2B_0/dff3B_6/Qb gnd! 2.1fF
C339 SubB_0/SR2B_0/dff3B_6/gate_2/Gin gnd! 16.9fF
C340 SubB_0/SR2B_0/dff3B_6/gate_2/Gout gnd! 4.4fF
C341 SubB_0/SR2B_0/dff3B_6/gate_1/Gin gnd! 17.3fF
C342 SubB_0/SR2B_0/dff3B_6/gate_3/Gin gnd! 17.4fF
C343 SubB_0/SR2B_0/dff3B_6/gate_3/Gout gnd! 4.4fF
C344 SubB_0/SR2B_0/dff3B_6/gate_0/S gnd! 26.8fF
C345 SubB_0/SR2B_0/dff3B_6/gate_2/S gnd! 33.8fF
C346 SubB_0/SR2B_0/dff3B_6/gate_1/S gnd! 27.4fF
C347 SubB_0/SR2B_0/dff3B_7/D gnd! 21.7fF
C348 SubB_0/SR2B_0/dff3B_7/inverter_7/out gnd! 11.5fF
C349 SubB_0/SR2B_0/dff3B_7/inverter_11/in gnd! 10.5fF
C350 SubB_0/SR2B_0/dff3B_7/gate_0/Gin gnd! 6.2fF
C351 SubB_0/SR2B_0/dff3B_7/Qb gnd! 2.1fF
C352 SubB_0/SR2B_0/dff3B_7/gate_2/Gin gnd! 16.9fF
C353 SubB_0/SR2B_0/dff3B_7/gate_2/Gout gnd! 4.4fF
C354 SubB_0/SR2B_0/dff3B_7/gate_1/Gin gnd! 17.3fF
C355 SubB_0/SR2B_0/dff3B_7/gate_3/Gin gnd! 17.4fF
C356 SubB_0/SR2B_0/dff3B_7/gate_3/Gout gnd! 4.4fF
C357 SubB_0/SR2B_0/dff3B_7/gate_0/S gnd! 26.8fF
C358 SubB_0/SR2B_0/dff3B_7/gate_2/S gnd! 33.8fF
C359 SubB_0/SR2B_0/dff3B_7/gate_1/S gnd! 27.4fF
C360 SubB_0/xor2_0/nand2_3/nand_in2 gnd! 28.1fF
C361 Cout gnd! 4.1fF
C362 SubB_0/xor2_0/nand2_4/nand_in2 gnd! 17.8fF
C363 SubB_0/xor2_0/nand2_4/nand_in1 gnd! 12.2fF
C364 SubB_0/dff3B_0/inverter_7/out gnd! 11.5fF
C365 SubB_0/dff3B_0/inverter_11/in gnd! 10.5fF
C366 SubB_0/dff3B_0/gate_0/Gin gnd! 6.2fF
C367 SubB_0/dff3B_0/Qb gnd! 2.1fF
C368 SubB_0/dff3B_0/gate_2/Gin gnd! 16.9fF
C369 SubB_0/dff3B_0/gate_2/Gout gnd! 4.4fF
C370 SubB_0/dff3B_0/gate_1/Gin gnd! 17.3fF
C371 SubB_0/dff3B_0/gate_3/Gin gnd! 17.4fF
C372 SubB_0/dff3B_0/gate_0/S gnd! 26.8fF
C373 SubB_0/dff3B_0/gate_2/S gnd! 33.8fF
C374 SubB_0/dff3B_0/gate_1/S gnd! 26.8fF
C375 SubB_0/SR2B_1/mux4x1_0/mux2x1_1/Smb gnd! 39.1fF
C376 SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Smb gnd! 22.7fF
C377 B0 gnd! 3.7fF
C378 SR2 gnd! 3.7fF
C379 SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Min1 gnd! 9.7fF
C380 SubB_0/SR2B_1/mux4x1_0/mux2x1_2/Min2 gnd! 12.2fF
C381 SubB_0/SR2B_1/mux4x1_1/mux2x1_1/Smb gnd! 39.1fF
C382 SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Smb gnd! 22.7fF
C383 B1 gnd! 3.7fF
C384 SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Min1 gnd! 9.7fF
C385 SubB_0/SR2B_1/mux4x1_1/mux2x1_2/Min2 gnd! 12.2fF
C386 SubB_0/SR2B_1/mux4x1_2/mux2x1_1/Smb gnd! 39.1fF
C387 SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Smb gnd! 22.7fF
C388 B2 gnd! 3.7fF
C389 SubB_0/SR2B_1/Q1 gnd! 146.9fF
C390 SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Min1 gnd! 9.7fF
C391 SubB_0/SR2B_1/mux4x1_2/mux2x1_2/Min2 gnd! 12.2fF
C392 SubB_0/SR2B_1/mux4x1_3/mux2x1_1/Smb gnd! 39.1fF
C393 SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Smb gnd! 22.7fF
C394 B3 gnd! 3.7fF
C395 SubB_0/SR2B_1/Q2 gnd! 134.6fF
C396 SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Min1 gnd! 9.7fF
C397 SubB_0/SR2B_1/mux4x1_3/mux2x1_2/Min2 gnd! 12.2fF
C398 SubB_0/SR2B_1/mux4x1_4/mux2x1_1/Smb gnd! 39.1fF
C399 SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Smb gnd! 22.7fF
C400 B4 gnd! 3.7fF
C401 SubB_0/SR2B_1/Q3 gnd! 146.9fF
C402 SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Min1 gnd! 9.7fF
C403 SubB_0/SR2B_1/mux4x1_4/mux2x1_2/Min2 gnd! 12.2fF
C404 SubB_0/SR2B_1/mux4x1_5/mux2x1_1/Smb gnd! 39.1fF
C405 SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Smb gnd! 22.7fF
C406 B5 gnd! 3.7fF
C407 SubB_0/SR2B_1/Q4 gnd! 134.6fF
C408 SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Min1 gnd! 9.7fF
C409 SubB_0/SR2B_1/mux4x1_5/mux2x1_2/Min2 gnd! 12.2fF
C410 SubB_0/SR2B_1/mux4x1_6/mux2x1_1/Smb gnd! 39.1fF
C411 SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Smb gnd! 22.7fF
C412 B6 gnd! 3.7fF
C413 SubB_0/SR2B_1/Q5 gnd! 118.7fF
C414 SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Min1 gnd! 9.7fF
C415 SubB_0/SR2B_1/mux4x1_6/mux2x1_2/Min2 gnd! 12.2fF
C416 SubB_0/SR2B_1/mux4x1_7/mux2x1_1/Smb gnd! 39.1fF
C417 SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Smb gnd! 22.7fF
C418 B7 gnd! 3.7fF
C419 SubB_0/SR2B_1/Q6 gnd! 134.6fF
C420 SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Min1 gnd! 9.7fF
C421 SubB_0/QB0 gnd! 299.6fF
C422 SubB_0/SR2B_1/mux4x1_7/mux2x1_2/Min2 gnd! 12.2fF
C423 SubB_0/SR2B_1/Q7 gnd! 115.7fF
C424 SubB_0/SR2B_1/dff3B_0/D gnd! 21.7fF
C425 SubB_0/SR2B_1/dff3B_0/inverter_7/out gnd! 11.5fF
C426 SubB_0/SR2B_1/dff3B_0/inverter_11/in gnd! 10.5fF
C427 SubB_0/SR2B_1/dff3B_0/gate_0/Gin gnd! 6.2fF
C428 SubB_0/SR2B_1/dff3B_0/Qb gnd! 2.1fF
C429 SubB_0/SR2B_1/dff3B_0/gate_2/Gin gnd! 16.9fF
C430 SubB_0/SR2B_1/dff3B_0/gate_2/Gout gnd! 4.4fF
C431 SubB_0/SR2B_1/dff3B_0/gate_1/Gin gnd! 17.3fF
C432 SubB_0/SR2B_1/dff3B_0/gate_3/Gin gnd! 17.4fF
C433 SubB_0/SR2B_1/dff3B_0/gate_3/Gout gnd! 4.4fF
C434 SubB_0/SR2B_1/dff3B_0/gate_0/S gnd! 26.8fF
C435 SubB_0/SR2B_1/dff3B_0/gate_2/S gnd! 33.8fF
C436 SubB_0/SR2B_1/dff3B_0/gate_1/S gnd! 27.4fF
C437 SubB_0/SR2B_1/dff3B_1/D gnd! 21.7fF
C438 SubB_0/SR2B_1/dff3B_1/inverter_7/out gnd! 11.5fF
C439 SubB_0/SR2B_1/dff3B_1/inverter_11/in gnd! 10.5fF
C440 SubB_0/SR2B_1/dff3B_1/gate_0/Gin gnd! 6.2fF
C441 SubB_0/SR2B_1/dff3B_1/Qb gnd! 2.1fF
C442 SubB_0/SR2B_1/dff3B_1/gate_2/Gin gnd! 16.9fF
C443 SubB_0/SR2B_1/dff3B_1/gate_2/Gout gnd! 4.4fF
C444 SubB_0/SR2B_1/dff3B_1/gate_1/Gin gnd! 17.3fF
C445 SubB_0/SR2B_1/dff3B_1/gate_3/Gin gnd! 17.4fF
C446 SubB_0/SR2B_1/dff3B_1/gate_3/Gout gnd! 4.4fF
C447 SubB_0/SR2B_1/dff3B_1/gate_0/S gnd! 26.8fF
C448 SubB_0/SR2B_1/dff3B_1/gate_2/S gnd! 33.8fF
C449 SubB_0/SR2B_1/dff3B_1/gate_1/S gnd! 27.4fF
C450 SubB_0/SR2B_1/dff3B_2/D gnd! 21.7fF
C451 SubB_0/SR2B_1/dff3B_2/inverter_7/out gnd! 11.5fF
C452 SubB_0/SR2B_1/dff3B_2/inverter_11/in gnd! 10.5fF
C453 SubB_0/SR2B_1/dff3B_2/gate_0/Gin gnd! 6.2fF
C454 SubB_0/SR2B_1/dff3B_2/Qb gnd! 2.1fF
C455 SubB_0/SR2B_1/dff3B_2/gate_2/Gin gnd! 16.9fF
C456 SubB_0/SR2B_1/dff3B_2/gate_2/Gout gnd! 4.4fF
C457 SubB_0/SR2B_1/dff3B_2/gate_1/Gin gnd! 17.3fF
C458 SubB_0/SR2B_1/dff3B_2/gate_3/Gin gnd! 17.4fF
C459 SubB_0/SR2B_1/dff3B_2/gate_3/Gout gnd! 4.4fF
C460 SubB_0/SR2B_1/dff3B_2/gate_0/S gnd! 26.8fF
C461 SubB_0/SR2B_1/dff3B_2/gate_2/S gnd! 33.8fF
C462 SubB_0/SR2B_1/dff3B_2/gate_1/S gnd! 27.4fF
C463 SubB_0/SR2B_1/dff3B_3/D gnd! 21.7fF
C464 SubB_0/SR2B_1/dff3B_3/inverter_7/out gnd! 11.5fF
C465 SubB_0/SR2B_1/dff3B_3/inverter_11/in gnd! 10.5fF
C466 SubB_0/SR2B_1/dff3B_3/gate_0/Gin gnd! 6.2fF
C467 SubB_0/SR2B_1/dff3B_3/Qb gnd! 2.1fF
C468 SubB_0/SR2B_1/dff3B_3/gate_2/Gin gnd! 16.9fF
C469 SubB_0/SR2B_1/dff3B_3/gate_2/Gout gnd! 4.4fF
C470 SubB_0/SR2B_1/dff3B_3/gate_1/Gin gnd! 17.3fF
C471 SubB_0/SR2B_1/dff3B_3/gate_3/Gin gnd! 17.4fF
C472 SubB_0/SR2B_1/dff3B_3/gate_3/Gout gnd! 4.4fF
C473 SubB_0/SR2B_1/dff3B_3/gate_0/S gnd! 26.8fF
C474 SubB_0/SR2B_1/dff3B_3/gate_2/S gnd! 33.8fF
C475 SubB_0/SR2B_1/dff3B_3/gate_1/S gnd! 27.4fF
C476 SubB_0/SR2B_1/dff3B_4/D gnd! 21.7fF
C477 SubB_0/SR2B_1/dff3B_4/inverter_7/out gnd! 11.5fF
C478 SubB_0/SR2B_1/dff3B_4/inverter_11/in gnd! 10.5fF
C479 SubB_0/SR2B_1/dff3B_4/gate_0/Gin gnd! 6.2fF
C480 SubB_0/SR2B_1/dff3B_4/Qb gnd! 2.1fF
C481 SubB_0/SR2B_1/dff3B_4/gate_2/Gin gnd! 16.9fF
C482 SubB_0/SR2B_1/dff3B_4/gate_2/Gout gnd! 4.4fF
C483 SubB_0/SR2B_1/dff3B_4/gate_1/Gin gnd! 17.3fF
C484 SubB_0/SR2B_1/dff3B_4/gate_3/Gin gnd! 17.4fF
C485 SubB_0/SR2B_1/dff3B_4/gate_3/Gout gnd! 4.4fF
C486 SubB_0/SR2B_1/dff3B_4/gate_0/S gnd! 26.8fF
C487 SubB_0/SR2B_1/dff3B_4/gate_2/S gnd! 33.8fF
C488 SubB_0/SR2B_1/dff3B_4/gate_1/S gnd! 27.4fF
C489 SubB_0/SR2B_1/dff3B_5/D gnd! 21.7fF
C490 SubB_0/SR2B_1/dff3B_5/inverter_7/out gnd! 11.5fF
C491 SubB_0/SR2B_1/dff3B_5/inverter_11/in gnd! 10.5fF
C492 SubB_0/SR2B_1/dff3B_5/gate_0/Gin gnd! 6.2fF
C493 SubB_0/SR2B_1/dff3B_5/Qb gnd! 2.1fF
C494 SubB_0/SR2B_1/dff3B_5/gate_2/Gin gnd! 16.9fF
C495 SubB_0/SR2B_1/dff3B_5/gate_2/Gout gnd! 4.4fF
C496 SubB_0/SR2B_1/dff3B_5/gate_1/Gin gnd! 17.3fF
C497 SubB_0/SR2B_1/dff3B_5/gate_3/Gin gnd! 17.4fF
C498 SubB_0/SR2B_1/dff3B_5/gate_3/Gout gnd! 4.4fF
C499 SubB_0/SR2B_1/dff3B_5/gate_0/S gnd! 26.8fF
C500 SubB_0/SR2B_1/dff3B_5/gate_2/S gnd! 33.8fF
C501 SubB_0/SR2B_1/dff3B_5/gate_1/S gnd! 27.4fF
C502 SubB_0/SR2B_1/dff3B_6/D gnd! 21.7fF
C503 SubB_0/SR2B_1/dff3B_6/inverter_7/out gnd! 11.5fF
C504 SubB_0/SR2B_1/dff3B_6/inverter_11/in gnd! 10.5fF
C505 SubB_0/SR2B_1/dff3B_6/gate_0/Gin gnd! 6.2fF
C506 SubB_0/SR2B_1/dff3B_6/Qb gnd! 2.1fF
C507 SubB_0/SR2B_1/dff3B_6/gate_2/Gin gnd! 16.9fF
C508 SubB_0/SR2B_1/dff3B_6/gate_2/Gout gnd! 4.4fF
C509 SubB_0/SR2B_1/dff3B_6/gate_1/Gin gnd! 17.3fF
C510 SubB_0/SR2B_1/dff3B_6/gate_3/Gin gnd! 17.4fF
C511 SubB_0/SR2B_1/dff3B_6/gate_3/Gout gnd! 4.4fF
C512 SubB_0/SR2B_1/dff3B_6/gate_0/S gnd! 26.8fF
C513 SubB_0/SR2B_1/dff3B_6/gate_2/S gnd! 33.8fF
C514 SubB_0/SR2B_1/dff3B_6/gate_1/S gnd! 27.4fF
C515 SubB_0/SR2B_1/dff3B_7/D gnd! 21.7fF
C516 SubB_0/SR2B_1/dff3B_7/inverter_7/out gnd! 11.5fF
C517 SubB_0/SR2B_1/dff3B_7/inverter_11/in gnd! 10.5fF
C518 SubB_0/SR2B_1/dff3B_7/gate_0/Gin gnd! 6.2fF
C519 SubB_0/SR2B_1/dff3B_7/Qb gnd! 2.1fF
C520 SubB_0/SR2B_1/dff3B_7/gate_2/Gin gnd! 16.9fF
C521 SubB_0/SR2B_1/dff3B_7/gate_2/Gout gnd! 4.4fF
C522 SubB_0/SR2B_1/dff3B_7/gate_1/Gin gnd! 17.3fF
C523 SubB_0/SR2B_1/dff3B_7/gate_3/Gin gnd! 17.4fF
C524 SubB_0/SR2B_1/dff3B_7/gate_3/Gout gnd! 4.4fF
C525 SubB_0/SR2B_1/dff3B_7/gate_0/S gnd! 26.8fF
C526 SubB_0/SR2B_1/dff3B_7/gate_2/S gnd! 33.8fF
C527 SubB_0/SR2B_1/dff3B_7/gate_1/S gnd! 27.4fF
C528 SubB_0/SR2B_2/mux4x1_0/mux2x1_1/Smb gnd! 39.1fF
C529 SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Smb gnd! 22.7fF
C530 D0 gnd! 3.7fF
C531 SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Min1 gnd! 9.7fF
C532 SubB_0/SR2B_2/mux4x1_0/mux2x1_2/Min2 gnd! 12.2fF
C533 SubB_0/SR2B_2/mux4x1_1/mux2x1_1/Smb gnd! 39.1fF
C534 SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Smb gnd! 22.7fF
C535 D1 gnd! 3.7fF
C536 SUM7 gnd! 89.6fF
C537 SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Min1 gnd! 9.7fF
C538 SubB_0/SR2B_2/mux4x1_1/mux2x1_2/Min2 gnd! 12.2fF
C539 SubB_0/SR2B_2/mux4x1_2/mux2x1_1/Smb gnd! 39.1fF
C540 SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Smb gnd! 22.7fF
C541 D2 gnd! 3.7fF
C542 SUM6 gnd! 146.9fF
C543 SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Min1 gnd! 9.7fF
C544 SubB_0/SR2B_2/mux4x1_2/mux2x1_2/Min2 gnd! 12.2fF
C545 SubB_0/SR2B_2/mux4x1_3/mux2x1_1/Smb gnd! 39.1fF
C546 SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Smb gnd! 22.7fF
C547 D3 gnd! 3.7fF
C548 SUM5 gnd! 134.6fF
C549 SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Min1 gnd! 9.7fF
C550 SubB_0/SR2B_2/mux4x1_3/mux2x1_2/Min2 gnd! 12.2fF
C551 SubB_0/SR2B_2/mux4x1_4/mux2x1_1/Smb gnd! 39.1fF
C552 SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Smb gnd! 22.7fF
C553 D4 gnd! 3.7fF
C554 SUM4 gnd! 146.9fF
C555 SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Min1 gnd! 9.7fF
C556 SubB_0/SR2B_2/mux4x1_4/mux2x1_2/Min2 gnd! 12.2fF
C557 SubB_0/SR2B_2/mux4x1_5/mux2x1_1/Smb gnd! 39.1fF
C558 SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Smb gnd! 22.7fF
C559 D5 gnd! 3.7fF
C560 SUM3 gnd! 134.6fF
C561 SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Min1 gnd! 9.7fF
C562 SubB_0/SR2B_2/mux4x1_5/mux2x1_2/Min2 gnd! 12.2fF
C563 SubB_0/SR2B_2/mux4x1_6/mux2x1_1/Smb gnd! 39.1fF
C564 SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Smb gnd! 22.7fF
C565 D6 gnd! 3.7fF
C566 SUM2 gnd! 118.7fF
C567 SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Min1 gnd! 9.7fF
C568 SubB_0/SR2B_2/mux4x1_6/mux2x1_2/Min2 gnd! 12.2fF
C569 SubB_0/SR2B_2/mux4x1_7/mux2x1_1/Smb gnd! 39.1fF
C570 nor2_0/out gnd! 496.1fF
C571 SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Smb gnd! 22.7fF
C572 D7 gnd! 3.7fF
C573 SUM1 gnd! 134.6fF
C574 SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Min1 gnd! 9.7fF
C575 SL gnd! 3.7fF
C576 SubB_0/SR2B_2/mux4x1_7/mux2x1_2/Min2 gnd! 12.2fF
C577 SUM0 gnd! 115.7fF
C578 SubB_0/SR2B_2/dff3B_0/D gnd! 21.7fF
C579 SubB_0/SR2B_2/dff3B_0/inverter_7/out gnd! 11.5fF
C580 SubB_0/SR2B_2/dff3B_0/inverter_11/in gnd! 10.5fF
C581 SubB_0/SR2B_2/dff3B_0/gate_0/Gin gnd! 6.2fF
C582 SubB_0/SR2B_2/dff3B_0/Qb gnd! 2.1fF
C583 SubB_0/SR2B_2/dff3B_0/gate_2/Gin gnd! 16.9fF
C584 SubB_0/SR2B_2/dff3B_0/gate_2/Gout gnd! 4.4fF
C585 SubB_0/SR2B_2/dff3B_0/gate_1/Gin gnd! 17.3fF
C586 SubB_0/SR2B_2/dff3B_0/gate_3/Gin gnd! 17.4fF
C587 SubB_0/SR2B_2/dff3B_0/gate_3/Gout gnd! 4.4fF
C588 SubB_0/SR2B_2/dff3B_0/gate_0/S gnd! 26.8fF
C589 SubB_0/SR2B_2/dff3B_0/gate_2/S gnd! 33.8fF
C590 SubB_0/SR2B_2/dff3B_0/gate_1/S gnd! 27.4fF
C591 SubB_0/SR2B_2/dff3B_1/D gnd! 21.7fF
C592 SubB_0/SR2B_2/dff3B_1/inverter_7/out gnd! 11.5fF
C593 SubB_0/SR2B_2/dff3B_1/inverter_11/in gnd! 10.5fF
C594 SubB_0/SR2B_2/dff3B_1/gate_0/Gin gnd! 6.2fF
C595 SubB_0/SR2B_2/dff3B_1/Qb gnd! 2.1fF
C596 SubB_0/SR2B_2/dff3B_1/gate_2/Gin gnd! 16.9fF
C597 SubB_0/SR2B_2/dff3B_1/gate_2/Gout gnd! 4.4fF
C598 SubB_0/SR2B_2/dff3B_1/gate_1/Gin gnd! 17.3fF
C599 SubB_0/SR2B_2/dff3B_1/gate_3/Gin gnd! 17.4fF
C600 SubB_0/SR2B_2/dff3B_1/gate_3/Gout gnd! 4.4fF
C601 SubB_0/SR2B_2/dff3B_1/gate_0/S gnd! 26.8fF
C602 SubB_0/SR2B_2/dff3B_1/gate_2/S gnd! 33.8fF
C603 SubB_0/SR2B_2/dff3B_1/gate_1/S gnd! 27.4fF
C604 SubB_0/SR2B_2/dff3B_2/D gnd! 21.7fF
C605 SubB_0/SR2B_2/dff3B_2/inverter_7/out gnd! 11.5fF
C606 SubB_0/SR2B_2/dff3B_2/inverter_11/in gnd! 10.5fF
C607 SubB_0/SR2B_2/dff3B_2/gate_0/Gin gnd! 6.2fF
C608 SubB_0/SR2B_2/dff3B_2/Qb gnd! 2.1fF
C609 SubB_0/SR2B_2/dff3B_2/gate_2/Gin gnd! 16.9fF
C610 SubB_0/SR2B_2/dff3B_2/gate_2/Gout gnd! 4.4fF
C611 SubB_0/SR2B_2/dff3B_2/gate_1/Gin gnd! 17.3fF
C612 SubB_0/SR2B_2/dff3B_2/gate_3/Gin gnd! 17.4fF
C613 SubB_0/SR2B_2/dff3B_2/gate_3/Gout gnd! 4.4fF
C614 SubB_0/SR2B_2/dff3B_2/gate_0/S gnd! 26.8fF
C615 SubB_0/SR2B_2/dff3B_2/gate_2/S gnd! 33.8fF
C616 SubB_0/SR2B_2/dff3B_2/gate_1/S gnd! 27.4fF
C617 SubB_0/SR2B_2/dff3B_3/D gnd! 21.7fF
C618 SubB_0/SR2B_2/dff3B_3/inverter_7/out gnd! 11.5fF
C619 SubB_0/SR2B_2/dff3B_3/inverter_11/in gnd! 10.5fF
C620 SubB_0/SR2B_2/dff3B_3/gate_0/Gin gnd! 6.2fF
C621 SubB_0/SR2B_2/dff3B_3/Qb gnd! 2.1fF
C622 SubB_0/SR2B_2/dff3B_3/gate_2/Gin gnd! 16.9fF
C623 SubB_0/SR2B_2/dff3B_3/gate_2/Gout gnd! 4.4fF
C624 SubB_0/SR2B_2/dff3B_3/gate_1/Gin gnd! 17.3fF
C625 SubB_0/SR2B_2/dff3B_3/gate_3/Gin gnd! 17.4fF
C626 SubB_0/SR2B_2/dff3B_3/gate_3/Gout gnd! 4.4fF
C627 SubB_0/SR2B_2/dff3B_3/gate_0/S gnd! 26.8fF
C628 SubB_0/SR2B_2/dff3B_3/gate_2/S gnd! 33.8fF
C629 SubB_0/SR2B_2/dff3B_3/gate_1/S gnd! 27.4fF
C630 SubB_0/SR2B_2/dff3B_4/D gnd! 21.7fF
C631 SubB_0/SR2B_2/dff3B_4/inverter_7/out gnd! 11.5fF
C632 SubB_0/SR2B_2/dff3B_4/inverter_11/in gnd! 10.5fF
C633 SubB_0/SR2B_2/dff3B_4/gate_0/Gin gnd! 6.2fF
C634 SubB_0/SR2B_2/dff3B_4/Qb gnd! 2.1fF
C635 SubB_0/SR2B_2/dff3B_4/gate_2/Gin gnd! 16.9fF
C636 SubB_0/SR2B_2/dff3B_4/gate_2/Gout gnd! 4.4fF
C637 SubB_0/SR2B_2/dff3B_4/gate_1/Gin gnd! 17.3fF
C638 SubB_0/SR2B_2/dff3B_4/gate_3/Gin gnd! 17.4fF
C639 SubB_0/SR2B_2/dff3B_4/gate_3/Gout gnd! 4.4fF
C640 SubB_0/SR2B_2/dff3B_4/gate_0/S gnd! 26.8fF
C641 SubB_0/SR2B_2/dff3B_4/gate_2/S gnd! 33.8fF
C642 SubB_0/SR2B_2/dff3B_4/gate_1/S gnd! 27.4fF
C643 SubB_0/SR2B_2/dff3B_5/D gnd! 21.7fF
C644 SubB_0/SR2B_2/dff3B_5/inverter_7/out gnd! 11.5fF
C645 SubB_0/SR2B_2/dff3B_5/inverter_11/in gnd! 10.5fF
C646 SubB_0/SR2B_2/dff3B_5/gate_0/Gin gnd! 6.2fF
C647 SubB_0/SR2B_2/dff3B_5/Qb gnd! 2.1fF
C648 SubB_0/SR2B_2/dff3B_5/gate_2/Gin gnd! 16.9fF
C649 SubB_0/SR2B_2/dff3B_5/gate_2/Gout gnd! 4.4fF
C650 SubB_0/SR2B_2/dff3B_5/gate_1/Gin gnd! 17.3fF
C651 SubB_0/SR2B_2/dff3B_5/gate_3/Gin gnd! 17.4fF
C652 SubB_0/SR2B_2/dff3B_5/gate_3/Gout gnd! 4.4fF
C653 SubB_0/SR2B_2/dff3B_5/gate_0/S gnd! 26.8fF
C654 SubB_0/SR2B_2/dff3B_5/gate_2/S gnd! 33.8fF
C655 SubB_0/SR2B_2/dff3B_5/gate_1/S gnd! 27.4fF
C656 SubB_0/SR2B_2/dff3B_6/D gnd! 21.7fF
C657 SubB_0/SR2B_2/dff3B_6/inverter_7/out gnd! 11.5fF
C658 SubB_0/SR2B_2/dff3B_6/inverter_11/in gnd! 10.5fF
C659 SubB_0/SR2B_2/dff3B_6/gate_0/Gin gnd! 6.2fF
C660 SubB_0/SR2B_2/dff3B_6/Qb gnd! 2.1fF
C661 SubB_0/SR2B_2/dff3B_6/gate_2/Gin gnd! 16.9fF
C662 SubB_0/SR2B_2/dff3B_6/gate_2/Gout gnd! 4.4fF
C663 SubB_0/SR2B_2/dff3B_6/gate_1/Gin gnd! 17.3fF
C664 SubB_0/SR2B_2/dff3B_6/gate_3/Gin gnd! 17.4fF
C665 SubB_0/SR2B_2/dff3B_6/gate_3/Gout gnd! 4.4fF
C666 SubB_0/SR2B_2/dff3B_6/gate_0/S gnd! 26.8fF
C667 SubB_0/SR2B_2/dff3B_6/gate_2/S gnd! 33.8fF
C668 SubB_0/SR2B_2/dff3B_6/gate_1/S gnd! 27.4fF
C669 SubB_0/SR2B_2/dff3B_7/D gnd! 21.7fF
C670 SubB_0/SR2B_2/dff3B_7/inverter_7/out gnd! 11.5fF
C671 SubB_0/SR2B_2/dff3B_7/inverter_11/in gnd! 10.5fF
C672 SubB_0/SR2B_2/dff3B_7/gate_0/Gin gnd! 6.2fF
C673 SubB_0/SR2B_2/dff3B_7/Qb gnd! 2.1fF
C674 SubB_0/SR2B_2/dff3B_7/gate_2/Gin gnd! 16.9fF
C675 SubB_0/SR2B_2/dff3B_7/gate_2/Gout gnd! 4.4fF
C676 SubB_0/SR2B_2/dff3B_7/gate_1/Gin gnd! 17.3fF
C677 SubB_0/SR2B_2/dff3B_7/gate_3/Gin gnd! 17.4fF
C678 SubB_0/SR2B_2/dff3B_7/gate_3/Gout gnd! 4.4fF
C679 SubB_0/SR2B_2/dff3B_7/gate_0/S gnd! 26.8fF
C680 SubB_0/SR2B_2/dff3B_7/gate_2/S gnd! 33.8fF
C681 SubB_0/SR2B_2/dff3B_7/gate_1/S gnd! 27.4fF

.include ../usc-spice

Vgnd1 GND 0 DC 0V
Vgnd2 gnd! 0 DC 0V
VVdd Vdd 0 DC 2.8V

Vin1 CLK 0 pulse(0 2.8 2ns 0.1ns 0.1ns 70ns 140ns)
Vin2 RST 0 pulse(0 2.8 120ns 0.1ns 0.1ns 140ns 2940ns)
Vin3 A0 0 pulse(2.8 2.8 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin4 A1 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin5 A2 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin6 A3 0 pulse(2.8 2.8 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin7 A4 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin8 A5 0 pulse(2.8 2.8 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin9 A6 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin10 A7 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin11 B0 0 pulse(2.8 2.8 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin12 B1 0 pulse(2.8 2.8 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin13 B2 0 pulse(2.8 2.8 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin14 B3 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin15 B4 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin16 B5 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin17 B6 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin18 B7 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin19 AbS 0 pulse(0 2.8 0ns 0.1ns 0.1ns 2940ns 5880ns)
Vin20 D0 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin21 D1 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin22 D2 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin23 D3 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin24 D4 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin25 D5 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin26 D6 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin27 D7 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin28 SR 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin29 SR2 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
Vin30 SL 0 pulse(0 0 0ns 0.1ns 0.1ns 5880ns 5880ns)
.tran 5ns 5880ns
.probe
.end
