magic
tech scmos
timestamp 1354203817
<< polysilicon >>
rect -11 308 -9 314
rect 30 309 32 321
rect 122 309 124 315
rect 163 309 165 321
rect 255 309 257 315
rect 296 309 298 321
rect 388 309 390 315
rect 429 309 431 321
rect 521 309 523 315
rect 562 309 564 321
rect 654 309 656 315
rect 695 309 697 321
rect 787 309 789 315
rect 828 309 830 321
rect 920 309 922 315
rect 961 309 963 321
rect 67 213 75 215
rect 200 213 208 215
rect 333 213 341 215
rect 466 213 474 215
rect 599 213 607 215
rect 732 213 740 215
rect 865 213 873 215
rect 998 213 1006 215
<< metal1 >>
rect 24 322 29 325
rect 33 322 162 325
rect 166 322 295 325
rect 299 322 428 325
rect 432 322 561 325
rect 565 322 694 325
rect 698 322 827 325
rect 831 322 960 325
rect -16 315 -12 318
rect -8 315 121 318
rect 125 315 254 318
rect 258 315 387 318
rect 391 315 520 318
rect 524 315 653 318
rect 657 315 786 318
rect 790 315 919 318
rect 90 309 219 312
rect 223 309 352 312
rect 356 309 485 312
rect 489 309 618 312
rect 622 309 751 312
rect 755 309 884 312
rect 888 309 1017 312
rect 26 302 120 305
rect 159 302 253 305
rect 292 302 386 305
rect 425 302 518 305
rect 558 302 652 305
rect 691 302 785 305
rect 824 302 918 305
rect 957 302 1029 305
rect -22 271 -18 274
rect 52 271 55 274
rect -22 230 -19 233
rect -22 -9 -19 218
rect 63 216 66 252
rect 79 239 82 278
rect 87 238 90 295
rect 95 238 98 302
rect 111 271 115 274
rect 185 271 188 274
rect 105 230 114 233
rect -6 58 -3 176
rect -6 55 3 58
rect 0 -3 3 55
rect 6 4 9 62
rect 105 29 108 230
rect 91 26 108 29
rect 14 10 17 22
rect 105 -3 108 26
rect 0 -6 108 -3
rect -22 -12 103 -9
rect 111 -15 114 218
rect 196 216 199 252
rect 212 239 215 278
rect 220 238 223 295
rect 228 238 231 302
rect 244 271 248 274
rect 318 271 321 274
rect 238 230 247 233
rect 127 58 130 176
rect 127 55 136 58
rect 133 -3 136 55
rect 139 4 142 62
rect 238 29 241 230
rect 224 26 241 29
rect 238 -3 241 26
rect 133 -6 241 -3
rect 133 -9 136 -6
rect 121 -12 136 -9
rect 244 -9 247 218
rect 329 216 332 252
rect 345 239 348 278
rect 353 238 356 295
rect 361 238 364 302
rect 377 271 381 274
rect 451 271 454 274
rect 371 230 380 233
rect 260 58 263 176
rect 260 55 269 58
rect 266 -2 269 55
rect 273 4 276 63
rect 371 29 374 230
rect 357 26 374 29
rect 371 -3 374 26
rect 269 -6 374 -3
rect 244 -12 369 -9
rect 377 -15 380 218
rect 462 216 465 252
rect 478 239 481 278
rect 486 238 489 295
rect 494 238 497 302
rect 510 271 514 274
rect 584 271 587 274
rect 504 230 513 233
rect 393 58 396 176
rect 393 55 402 58
rect 399 -3 402 55
rect 405 4 408 63
rect 504 29 507 230
rect 490 26 507 29
rect 504 -3 507 26
rect 399 -6 507 -3
rect 399 -9 402 -6
rect 387 -12 402 -9
rect 510 -9 513 218
rect 595 216 598 252
rect 611 239 614 278
rect 619 238 622 295
rect 627 238 630 302
rect 643 271 647 274
rect 717 271 720 274
rect 637 230 646 233
rect 526 58 529 176
rect 526 55 535 58
rect 532 -2 535 55
rect 539 4 542 62
rect 637 29 640 230
rect 623 26 640 29
rect 637 -3 640 26
rect 535 -6 640 -3
rect 510 -12 635 -9
rect 643 -15 646 218
rect 728 216 731 252
rect 744 239 747 278
rect 752 238 755 295
rect 760 238 763 302
rect 776 271 780 274
rect 850 271 853 274
rect 770 230 779 233
rect 659 58 662 176
rect 659 55 668 58
rect 665 -3 668 55
rect 671 4 674 62
rect 770 29 773 230
rect 756 26 773 29
rect 770 -3 773 26
rect 665 -6 773 -3
rect 665 -9 668 -6
rect 653 -12 668 -9
rect 776 -9 779 218
rect 861 216 864 252
rect 877 239 880 278
rect 885 238 888 295
rect 893 238 896 302
rect 909 271 913 274
rect 983 271 986 274
rect 903 230 912 233
rect 792 58 795 176
rect 792 55 801 58
rect 798 -2 801 55
rect 805 6 808 64
rect 903 29 906 230
rect 909 215 912 218
rect 994 216 997 252
rect 1010 239 1013 278
rect 1018 238 1021 295
rect 1026 238 1029 302
rect 925 58 928 176
rect 925 55 934 58
rect 889 26 906 29
rect 903 -3 906 26
rect 801 -6 906 -3
rect 931 -3 934 55
rect 937 4 940 62
rect 1022 26 1039 29
rect 1036 -3 1039 26
rect 931 -6 1039 -3
rect 931 -9 934 -6
rect 776 -12 934 -9
rect 111 -18 265 -15
rect 377 -18 531 -15
rect 643 -18 797 -15
rect 7 -22 10 -19
rect 7 -25 139 -22
rect 143 -25 273 -22
rect 277 -25 405 -22
rect 409 -25 539 -22
rect 543 -25 671 -22
rect 675 -24 805 -22
rect 809 -24 937 -22
rect 675 -25 940 -24
rect 17 -31 147 -28
rect 151 -31 281 -28
rect 285 -31 414 -28
rect 418 -31 547 -28
rect 551 -31 679 -28
rect 683 -31 813 -28
rect 817 -31 945 -28
<< metal2 >>
rect 87 299 90 308
rect 220 299 223 308
rect 353 299 356 308
rect 486 299 489 308
rect 619 299 622 308
rect 752 299 755 308
rect 885 299 888 308
rect 1018 299 1021 308
rect 3 279 78 282
rect 136 279 211 282
rect 269 279 344 282
rect 402 279 477 282
rect 535 279 610 282
rect 667 279 743 282
rect 800 279 876 282
rect 933 279 1009 282
rect 13 26 16 86
rect 147 15 150 87
rect 280 15 283 87
rect 413 15 416 87
rect 546 15 549 87
rect 678 15 681 87
rect 812 15 815 87
rect 147 12 151 15
rect 280 12 284 15
rect 413 12 417 15
rect 546 12 550 15
rect 678 12 682 15
rect 812 12 816 15
rect 6 -15 9 0
rect 14 -28 17 6
rect 107 -12 117 -9
rect 139 -21 142 0
rect 148 -28 151 12
rect 266 -15 269 -6
rect 273 -21 276 0
rect 281 -28 284 12
rect 373 -12 383 -9
rect 405 -21 408 0
rect 414 -28 417 12
rect 532 -15 535 -6
rect 539 -21 542 0
rect 547 -28 550 12
rect 639 -12 649 -9
rect 671 -21 674 0
rect 679 -28 682 12
rect 798 -15 801 -6
rect 805 -20 808 2
rect 813 -28 816 12
rect 937 -20 940 0
rect 945 -28 948 87
<< polycontact >>
rect 29 321 33 325
rect 162 321 166 325
rect 295 321 299 325
rect 428 321 432 325
rect 561 321 565 325
rect 694 321 698 325
rect 827 321 831 325
rect 960 321 964 325
rect -12 314 -8 318
rect 121 315 125 319
rect 254 315 258 319
rect 387 315 391 319
rect 520 315 524 319
rect 653 315 657 319
rect 786 315 790 319
rect 919 315 923 319
rect 86 234 90 238
rect 219 234 223 238
rect 352 234 356 238
rect 485 234 489 238
rect 618 234 622 238
rect 751 234 755 238
rect 884 234 888 238
rect 1017 234 1021 238
rect 63 212 67 216
rect 196 212 200 216
rect 329 212 333 216
rect 462 212 466 216
rect 595 212 599 216
rect 728 212 732 216
rect 861 212 865 216
rect 994 212 998 216
<< m2contact >>
rect 86 308 90 312
rect 219 308 223 312
rect 352 308 356 312
rect 485 308 489 312
rect 618 308 622 312
rect 751 308 755 312
rect 884 308 888 312
rect 1017 308 1021 312
rect 86 295 90 299
rect 78 278 82 282
rect 219 295 223 299
rect 211 278 215 282
rect 13 22 17 26
rect 14 6 18 10
rect 6 0 10 4
rect 103 -13 107 -9
rect 352 295 356 299
rect 344 278 348 282
rect 139 0 143 4
rect 117 -12 121 -8
rect 485 295 489 299
rect 477 278 481 282
rect 273 0 277 4
rect 265 -6 269 -2
rect 369 -13 373 -9
rect 618 295 622 299
rect 610 278 614 282
rect 405 0 409 4
rect 383 -12 387 -8
rect 751 295 755 299
rect 743 278 747 282
rect 539 0 543 4
rect 531 -6 535 -2
rect 635 -13 639 -9
rect 884 295 888 299
rect 876 278 880 282
rect 671 0 675 4
rect 649 -12 653 -8
rect 1017 295 1021 299
rect 1009 278 1013 282
rect 804 2 808 6
rect 797 -6 801 -2
rect 937 0 941 4
rect 6 -19 10 -15
rect 265 -19 269 -15
rect 531 -19 535 -15
rect 797 -19 801 -15
rect 139 -25 143 -21
rect 273 -25 277 -21
rect 405 -25 409 -21
rect 539 -25 543 -21
rect 671 -25 675 -21
rect 805 -24 809 -20
rect 937 -24 941 -20
rect 13 -32 17 -28
rect 147 -32 151 -28
rect 281 -32 285 -28
rect 414 -32 418 -28
rect 547 -32 551 -28
rect 679 -32 683 -28
rect 813 -32 817 -28
rect 945 -32 949 -28
use mux4x1 mux4x1_0
timestamp 1353620947
transform 1 0 -14 0 1 229
box -8 -56 80 81
use mux4x1 mux4x1_1
timestamp 1353620947
transform 1 0 119 0 1 229
box -8 -56 80 81
use mux4x1 mux4x1_2
timestamp 1353620947
transform 1 0 252 0 1 229
box -8 -56 80 81
use mux4x1 mux4x1_3
timestamp 1353620947
transform 1 0 385 0 1 229
box -8 -56 80 81
use mux4x1 mux4x1_4
timestamp 1353620947
transform 1 0 518 0 1 229
box -8 -56 80 81
use mux4x1 mux4x1_5
timestamp 1353620947
transform 1 0 651 0 1 229
box -8 -56 80 81
use mux4x1 mux4x1_6
timestamp 1353620947
transform 1 0 784 0 1 229
box -8 -56 80 81
use mux4x1 mux4x1_7
timestamp 1353620947
transform 1 0 917 0 1 229
box -8 -56 80 81
use dff3B dff3B_0
timestamp 1354117195
transform 0 1 72 -1 0 130
box -110 -72 130 37
use dff3B dff3B_1
timestamp 1354117195
transform 0 1 205 -1 0 130
box -110 -72 130 37
use dff3B dff3B_2
timestamp 1354117195
transform 0 1 338 -1 0 130
box -110 -72 130 37
use dff3B dff3B_3
timestamp 1354117195
transform 0 1 471 -1 0 130
box -110 -72 130 37
use dff3B dff3B_4
timestamp 1354117195
transform 0 1 604 -1 0 130
box -110 -72 130 37
use dff3B dff3B_5
timestamp 1354117195
transform 0 1 737 -1 0 130
box -110 -72 130 37
use dff3B dff3B_6
timestamp 1354117195
transform 0 1 870 -1 0 130
box -110 -72 130 37
use dff3B dff3B_7
timestamp 1354117195
transform 0 1 1003 -1 0 130
box -110 -72 130 37
<< labels >>
rlabel metal1 -14 316 -14 316 1 S1
rlabel metal1 26 323 26 323 5 S0
rlabel metal1 60 303 60 303 1 Vdd!
rlabel metal1 -20 273 -20 273 3 IN0
rlabel metal1 -21 232 -21 232 3 SR
rlabel metal1 113 273 113 273 1 IN1
rlabel metal1 246 273 246 273 1 IN2
rlabel metal1 380 273 380 273 1 IN3
rlabel metal1 512 273 512 273 1 IN4
rlabel metal1 645 273 645 273 1 IN5
rlabel metal1 778 273 778 273 1 IN6
rlabel metal1 911 273 911 273 1 IN7
rlabel metal1 8 -24 8 -24 1 CLK
rlabel metal1 27 -30 27 -30 1 GND!
rlabel metal1 97 310 97 310 1 CLR
rlabel metal1 106 27 106 27 1 Q0
rlabel metal1 240 27 240 27 1 Q1
rlabel metal1 372 27 372 27 1 Q2
rlabel metal1 505 27 505 27 1 Q3
rlabel metal1 638 27 638 27 1 Q4
rlabel metal1 771 27 771 27 1 Q5
rlabel metal1 904 27 904 27 1 Q6
rlabel metal1 1038 27 1038 27 7 Q7
rlabel metal1 911 217 911 217 1 SL
<< end >>
