magic
tech scmos
timestamp 1357664372
<< polysilicon >>
rect 212 1156 214 1159
rect 531 1157 533 1168
rect 51 879 54 881
rect 212 659 214 668
rect 236 659 238 668
<< metal1 >>
rect 147 1477 155 1480
rect 124 1461 127 1467
rect 65 1458 69 1461
rect 164 1456 168 1460
rect 1110 1457 1142 1460
rect 207 1161 210 1171
rect 241 1171 244 1189
rect 241 1168 266 1171
rect 55 1132 58 1159
rect 207 1158 228 1161
rect 207 1153 210 1158
rect 225 1153 228 1158
rect 218 1142 227 1145
rect 236 1141 250 1144
rect 247 1137 250 1141
rect 257 1137 260 1144
rect 207 1132 210 1137
rect 225 1132 228 1136
rect 247 1134 260 1137
rect 55 1129 228 1132
rect 236 996 239 1112
rect 48 993 239 996
rect 48 883 51 993
rect 257 737 260 1134
rect 263 1067 266 1168
rect 289 1109 292 1131
rect 369 1109 372 1125
rect 406 1102 409 1128
rect 418 1127 436 1130
rect 450 1127 457 1130
rect 418 1103 421 1127
rect 270 1099 409 1102
rect 270 1087 273 1099
rect 443 1096 446 1124
rect 454 1103 457 1127
rect 477 1124 480 1129
rect 529 1116 532 1153
rect 472 1113 532 1116
rect 276 1093 446 1096
rect 276 1079 279 1093
rect 293 1086 296 1089
rect 1331 1062 1334 1091
rect 413 1035 418 1038
rect 546 1035 551 1038
rect 679 1035 684 1038
rect 812 1035 817 1038
rect 945 1035 950 1038
rect 1078 1035 1083 1038
rect 1211 1035 1216 1038
rect 283 1032 286 1035
rect 283 991 286 994
rect 1347 733 1350 1021
rect 276 694 279 698
rect 65 683 68 687
rect 242 687 245 690
rect 238 684 245 687
rect 201 673 204 679
rect 218 677 225 679
rect 218 676 228 677
rect 201 670 211 673
rect 207 666 210 670
rect 223 666 226 671
rect 239 666 242 671
rect 282 666 285 671
rect 412 669 417 672
rect 545 669 553 672
rect 678 669 685 672
rect 811 669 816 672
rect 944 669 950 672
rect 1077 669 1084 672
rect 1210 669 1217 672
rect 207 663 242 666
rect 216 655 235 658
rect 235 628 238 655
rect 186 625 238 628
rect 282 625 285 630
rect 24 579 27 582
rect 282 300 285 304
rect 415 300 418 306
rect 548 300 551 306
rect 681 300 684 306
rect 814 300 817 306
rect 947 300 950 306
rect 1080 300 1083 306
rect 1213 300 1216 306
rect 1213 244 1216 250
rect 409 58 412 61
rect 542 58 545 61
rect 675 58 678 61
rect 808 58 811 61
rect 941 58 944 61
rect 1074 58 1077 61
rect 1207 58 1210 61
rect 1340 58 1343 61
<< metal2 >>
rect 55 1163 58 1297
rect 138 1175 141 1214
rect 1126 1213 1142 1216
rect 156 1206 244 1209
rect 241 1193 244 1206
rect 138 1172 206 1175
rect 257 1148 260 1199
rect 226 1120 476 1123
rect 226 702 229 1120
rect 240 1113 468 1116
rect 289 1090 292 1105
rect 369 1091 372 1105
rect 411 1099 417 1102
rect 445 1100 454 1103
rect 369 1088 403 1091
rect 400 1083 403 1088
rect 411 1069 414 1099
rect 445 1044 448 1100
rect 1347 1025 1350 1091
rect 226 699 276 702
rect 246 691 269 694
rect 211 685 223 688
rect 207 655 210 685
rect 235 655 239 659
<< polycontact >>
rect 529 1153 533 1157
rect 227 1142 231 1146
rect 47 879 51 883
rect 225 677 229 681
rect 212 655 216 659
rect 235 655 239 659
<< m2contact >>
rect 152 1206 156 1210
rect 256 1199 260 1203
rect 241 1189 245 1193
rect 206 1171 210 1175
rect 55 1159 59 1163
rect 256 1144 260 1148
rect 236 1112 240 1116
rect 289 1105 293 1109
rect 368 1105 372 1109
rect 417 1099 421 1103
rect 476 1120 480 1124
rect 468 1112 472 1116
rect 454 1099 458 1103
rect 289 1086 293 1090
rect 400 1079 404 1083
rect 410 1065 414 1069
rect 1346 1021 1350 1025
rect 276 698 280 702
rect 242 690 246 694
rect 269 690 273 694
rect 207 685 211 689
rect 223 685 227 689
use inverter inverter_2
timestamp 1351319193
transform 1 0 212 0 1 1142
box -5 -10 7 15
use inverter inverter_1
timestamp 1351319193
transform 1 0 230 0 1 1142
box -5 -10 7 15
use fsm fsm_0
timestamp 1354710338
transform 1 0 156 0 1 1200
box -159 -79 983 290
use inverter inverter_0
timestamp 1351319193
transform 1 0 212 0 1 676
box -5 -10 7 15
use nor2 nor2_0
timestamp 1351504687
transform 1 0 267 0 1 677
box -44 -11 -24 15
use SubB SubB_0
timestamp 1357465246
transform 1 0 283 0 1 732
box -283 -732 1074 357
<< labels >>
rlabel metal1 66 684 66 684 1 AbS
rlabel metal1 26 580 26 580 1 Cout
rlabel metal1 284 992 284 992 1 SR
rlabel metal1 285 1034 285 1034 1 A0
rlabel metal1 1214 1036 1214 1036 1 A7
rlabel metal1 1080 1036 1080 1036 1 A6
rlabel metal1 947 1037 947 1037 1 A5
rlabel metal1 814 1036 814 1036 1 A4
rlabel metal1 681 1037 681 1037 1 A3
rlabel metal1 547 1037 547 1037 1 A2
rlabel metal1 414 1037 414 1037 1 A1
rlabel metal1 283 667 283 667 1 B0
rlabel metal1 283 626 283 626 1 SR2
rlabel metal1 415 670 415 670 1 B1
rlabel metal1 548 670 548 670 1 B2
rlabel metal1 681 671 681 671 1 B3
rlabel metal1 814 670 814 670 1 B4
rlabel metal1 947 670 947 670 1 B5
rlabel metal1 1080 670 1080 670 1 B6
rlabel metal1 1213 670 1213 670 1 B7
rlabel metal1 283 302 283 302 1 D0
rlabel metal1 1215 302 1215 302 1 D7
rlabel metal1 1081 302 1081 302 1 D6
rlabel metal1 948 302 948 302 1 D5
rlabel metal1 816 302 816 302 1 D4
rlabel metal1 682 302 682 302 1 D3
rlabel metal1 549 302 549 302 1 D2
rlabel metal1 416 302 416 302 1 D1
rlabel metal1 1215 246 1215 246 1 SL
rlabel metal1 1341 59 1341 59 1 SUM0
rlabel metal1 1209 59 1209 59 1 SUM1
rlabel metal1 1076 59 1076 59 1 SUM2
rlabel metal1 943 59 943 59 1 SUM3
rlabel metal1 810 59 810 59 1 SUM4
rlabel metal1 677 59 677 59 1 SUM5
rlabel metal1 543 59 543 59 1 SUM6
rlabel metal1 411 59 411 59 1 SUM7
rlabel metal1 150 1478 150 1478 1 RST
rlabel metal1 290 1125 290 1125 1 SA0
rlabel metal1 371 1118 371 1118 1 SA1
rlabel metal1 407 1118 407 1118 1 SB0
rlabel metal1 444 1117 444 1117 1 SB1
rlabel metal1 478 1125 478 1125 1 SS0
rlabel metal1 125 1465 125 1465 1 GND!
rlabel metal1 66 1460 66 1460 1 Vdd!
rlabel polysilicon 213 1158 213 1158 1 CLK
<< end >>
