* SPICE3 file created from gate.ext - technology: scmos

M1000 Gout S Gin Vdd pfet w=6u l=2u
+ ad=49p pd=30u as=49p ps=30u 
M1001 Gout Sb Gin Gnd nfet w=3u l=2u
+ ad=28p pd=24u as=28p ps=24u 
C0 Sb gnd! 2.1fF
C1 S gnd! 2.1fF

.include ../usc-spice

Vgnd1 GND 0 DC 0V
Vgnd2 gnd! 0 DC 0V
VVdd Vdd 0 DC 2.8V

Vin1 S 0 pulse(2.8 0 0ns 0.1ns 0.1ns 5ns 10ns)
Vin2 Sb 0 pulse(0 2.8 0ns 0.1ns 0.1ns 5ns 10ns)
Vin3 Gin 0 pulse(0 2.8 0ns 0.1ns 0.1ns 10ns 20ns)
.tran 5ns 40ns
.probe
.end
