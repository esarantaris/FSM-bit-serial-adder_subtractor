magic
tech scmos
timestamp 1353094667
<< polysilicon >>
rect -1 17 1 20
rect -1 8 1 11
rect -1 1 1 4
rect -1 -5 1 -2
<< ndiffusion >>
rect -5 -2 -1 1
rect 1 -2 5 1
<< pdiffusion >>
rect -5 14 -1 17
rect -8 11 -1 14
rect 1 14 5 17
rect 1 11 8 14
<< metal1 >>
rect -8 1 -5 14
rect 5 1 8 14
<< ntransistor >>
rect -1 -2 1 1
<< ptransistor >>
rect -1 11 1 17
<< ndcontact >>
rect -9 -3 -5 1
rect 5 -3 9 1
<< pdcontact >>
rect -9 14 -5 18
rect 5 14 9 18
<< labels >>
rlabel polysilicon 0 19 0 19 5 S
rlabel polysilicon 0 -4 0 -4 1 Sb
rlabel metal1 -7 6 -7 6 3 Gin
rlabel metal1 7 6 7 6 7 Gout
<< end >>
