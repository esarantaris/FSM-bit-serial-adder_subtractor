magic
tech scmos
timestamp 1352389694
<< polysilicon >>
rect -36 18 -34 29
rect -28 22 -26 29
rect -28 20 3 22
rect -28 18 -26 20
rect 1 18 3 20
rect -36 -21 -34 -14
rect -20 -19 -18 -2
rect -32 -21 -18 -19
rect -3 -18 8 -16
rect -3 -21 -1 -18
<< metal1 >>
rect -41 23 21 26
rect -41 14 -38 23
rect -24 14 -21 23
rect -11 14 -8 23
rect 5 14 8 23
rect -25 -2 -20 1
rect -16 -2 -10 1
rect 4 -2 12 1
rect -40 -16 -37 -13
rect -11 -16 -8 -13
rect 9 -14 12 -2
rect -47 -19 -8 -16
rect -47 -62 -44 -19
rect -40 -22 -37 -19
rect -11 -22 -8 -19
rect -25 -38 -10 -35
rect 4 -38 11 -35
rect -40 -55 -37 -49
rect -24 -55 -21 -49
rect -11 -55 -8 -49
rect 5 -55 8 -49
rect 18 -55 21 23
rect -40 -58 21 -55
<< polycontact >>
rect -20 -2 -16 2
rect -10 -2 -6 2
rect 8 -18 12 -14
rect -10 -39 -6 -35
use nand2 nand2_1
timestamp 1288918752
transform 1 0 3 0 1 -6
box -44 -8 -24 24
use nand2 nand2_2
timestamp 1288918752
transform 1 0 32 0 1 -6
box -44 -8 -24 24
use nand2 nand2_3
timestamp 1288918752
transform 1 0 3 0 -1 -29
box -44 -8 -24 24
use nand2 nand2_4
timestamp 1288918752
transform 1 0 32 0 -1 -29
box -44 -8 -24 24
<< labels >>
rlabel polysilicon -27 27 -27 27 1 xor_in2
rlabel metal1 19 -17 19 -17 1 Vdd!
rlabel metal1 -46 -60 -46 -60 1 GND!
rlabel metal1 10 -37 10 -37 1 xor_out
rlabel polysilicon -35 27 -35 27 5 xor_in1
<< end >>
