magic
tech scmos
timestamp 1354114587
<< polysilicon >>
rect 11 129 13 132
rect 19 129 21 132
rect 11 91 13 97
rect 15 93 17 97
rect 15 91 21 93
rect 61 24 73 26
<< metal1 >>
rect 65 131 68 132
rect 6 128 68 131
rect 6 125 9 128
rect 23 125 26 128
rect 30 125 33 128
rect 22 112 32 115
rect 42 112 52 115
rect 6 95 9 98
rect 30 95 33 105
rect 0 92 33 95
rect 0 0 3 92
rect 65 88 68 128
<< polycontact >>
rect 32 112 36 116
rect 57 23 61 27
use nand2 nand2_0
timestamp 1288918752
transform 1 0 50 0 1 105
box -44 -8 -24 24
use not1 not1_0
timestamp 1352402877
transform 1 0 35 0 1 112
box -5 -10 7 15
use xor2 xor2_0
timestamp 1352389694
transform 1 0 47 0 1 62
box -47 -62 21 29
<< labels >>
rlabel polysilicon 12 131 12 131 5 ha_in1
rlabel polysilicon 20 131 20 131 5 ha_in2
rlabel polysilicon 72 25 72 25 7 ha_sum
rlabel metal1 51 113 51 113 7 ha_cout
rlabel metal1 66 128 66 128 5 Vdd!
rlabel metal1 2 94 2 94 3 GND!
<< end >>
